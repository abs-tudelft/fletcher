tb.hm_put_byte(.addr(0), .d(8'h00));
tb.hm_put_byte(.addr(1), .d(8'h00));
tb.hm_put_byte(.addr(2), .d(8'h00));
tb.hm_put_byte(.addr(3), .d(8'h00));
tb.hm_put_byte(.addr(4), .d(8'h08));
tb.hm_put_byte(.addr(5), .d(8'h00));
tb.hm_put_byte(.addr(6), .d(8'h00));
tb.hm_put_byte(.addr(7), .d(8'h00));
tb.hm_put_byte(.addr(8), .d(8'h10));
tb.hm_put_byte(.addr(9), .d(8'h00));
tb.hm_put_byte(.addr(10), .d(8'h00));
tb.hm_put_byte(.addr(11), .d(8'h00));
tb.hm_put_byte(.addr(12), .d(8'h18));
tb.hm_put_byte(.addr(13), .d(8'h00));
tb.hm_put_byte(.addr(14), .d(8'h00));
tb.hm_put_byte(.addr(15), .d(8'h00));
tb.hm_put_byte(.addr(16), .d(8'h20));
tb.hm_put_byte(.addr(17), .d(8'h00));
tb.hm_put_byte(.addr(18), .d(8'h00));
tb.hm_put_byte(.addr(19), .d(8'h00));
tb.hm_put_byte(.addr(20), .d(8'h28));
tb.hm_put_byte(.addr(21), .d(8'h00));
tb.hm_put_byte(.addr(22), .d(8'h00));
tb.hm_put_byte(.addr(23), .d(8'h00));
tb.hm_put_byte(.addr(24), .d(8'h00));
tb.hm_put_byte(.addr(25), .d(8'h00));
tb.hm_put_byte(.addr(26), .d(8'h00));
tb.hm_put_byte(.addr(27), .d(8'h00));
tb.hm_put_byte(.addr(28), .d(8'h00));
tb.hm_put_byte(.addr(29), .d(8'h00));
tb.hm_put_byte(.addr(30), .d(8'h00));
tb.hm_put_byte(.addr(31), .d(8'h00));
tb.hm_put_byte(.addr(32), .d(8'h00));
tb.hm_put_byte(.addr(33), .d(8'h00));
tb.hm_put_byte(.addr(34), .d(8'h00));
tb.hm_put_byte(.addr(35), .d(8'h00));
tb.hm_put_byte(.addr(36), .d(8'h00));
tb.hm_put_byte(.addr(37), .d(8'h00));
tb.hm_put_byte(.addr(38), .d(8'h00));
tb.hm_put_byte(.addr(39), .d(8'h00));
tb.hm_put_byte(.addr(40), .d(8'h00));
tb.hm_put_byte(.addr(41), .d(8'h00));
tb.hm_put_byte(.addr(42), .d(8'h00));
tb.hm_put_byte(.addr(43), .d(8'h00));
tb.hm_put_byte(.addr(44), .d(8'h00));
tb.hm_put_byte(.addr(45), .d(8'h00));
tb.hm_put_byte(.addr(46), .d(8'h00));
tb.hm_put_byte(.addr(47), .d(8'h00));
tb.hm_put_byte(.addr(48), .d(8'h00));
tb.hm_put_byte(.addr(49), .d(8'h00));
tb.hm_put_byte(.addr(50), .d(8'h00));
tb.hm_put_byte(.addr(51), .d(8'h00));
tb.hm_put_byte(.addr(52), .d(8'h00));
tb.hm_put_byte(.addr(53), .d(8'h00));
tb.hm_put_byte(.addr(54), .d(8'h00));
tb.hm_put_byte(.addr(55), .d(8'h00));
tb.hm_put_byte(.addr(56), .d(8'h00));
tb.hm_put_byte(.addr(57), .d(8'h00));
tb.hm_put_byte(.addr(58), .d(8'h00));
tb.hm_put_byte(.addr(59), .d(8'h00));
tb.hm_put_byte(.addr(60), .d(8'h00));
tb.hm_put_byte(.addr(61), .d(8'h00));
tb.hm_put_byte(.addr(62), .d(8'h00));
tb.hm_put_byte(.addr(63), .d(8'h00));
tb.hm_put_byte(.addr(64), .d(8'h0C));
tb.hm_put_byte(.addr(65), .d(8'h00));
tb.hm_put_byte(.addr(66), .d(8'h00));
tb.hm_put_byte(.addr(67), .d(8'h00));
tb.hm_put_byte(.addr(68), .d(8'h00));
tb.hm_put_byte(.addr(69), .d(8'h00));
tb.hm_put_byte(.addr(70), .d(8'h00));
tb.hm_put_byte(.addr(71), .d(8'h00));
tb.hm_put_byte(.addr(72), .d(8'h06));
tb.hm_put_byte(.addr(73), .d(8'h00));
tb.hm_put_byte(.addr(74), .d(8'h00));
tb.hm_put_byte(.addr(75), .d(8'h00));
tb.hm_put_byte(.addr(76), .d(8'h00));
tb.hm_put_byte(.addr(77), .d(8'h00));
tb.hm_put_byte(.addr(78), .d(8'h00));
tb.hm_put_byte(.addr(79), .d(8'h00));
tb.hm_put_byte(.addr(80), .d(8'h6E));
tb.hm_put_byte(.addr(81), .d(8'h00));
tb.hm_put_byte(.addr(82), .d(8'h00));
tb.hm_put_byte(.addr(83), .d(8'h00));
tb.hm_put_byte(.addr(84), .d(8'h00));
tb.hm_put_byte(.addr(85), .d(8'h00));
tb.hm_put_byte(.addr(86), .d(8'h00));
tb.hm_put_byte(.addr(87), .d(8'h00));
tb.hm_put_byte(.addr(88), .d(8'h78));
tb.hm_put_byte(.addr(89), .d(8'h00));
tb.hm_put_byte(.addr(90), .d(8'h00));
tb.hm_put_byte(.addr(91), .d(8'h00));
tb.hm_put_byte(.addr(92), .d(8'h00));
tb.hm_put_byte(.addr(93), .d(8'h00));
tb.hm_put_byte(.addr(94), .d(8'h00));
tb.hm_put_byte(.addr(95), .d(8'h00));
tb.hm_put_byte(.addr(96), .d(8'h82));
tb.hm_put_byte(.addr(97), .d(8'h00));
tb.hm_put_byte(.addr(98), .d(8'h00));
tb.hm_put_byte(.addr(99), .d(8'h00));
tb.hm_put_byte(.addr(100), .d(8'h00));
tb.hm_put_byte(.addr(101), .d(8'h00));
tb.hm_put_byte(.addr(102), .d(8'h00));
tb.hm_put_byte(.addr(103), .d(8'h00));
tb.hm_put_byte(.addr(104), .d(8'h8C));
tb.hm_put_byte(.addr(105), .d(8'h00));
tb.hm_put_byte(.addr(106), .d(8'h00));
tb.hm_put_byte(.addr(107), .d(8'h00));
tb.hm_put_byte(.addr(108), .d(8'h00));
tb.hm_put_byte(.addr(109), .d(8'h00));
tb.hm_put_byte(.addr(110), .d(8'h00));
tb.hm_put_byte(.addr(111), .d(8'h00));
tb.hm_put_byte(.addr(112), .d(8'h96));
tb.hm_put_byte(.addr(113), .d(8'h00));
tb.hm_put_byte(.addr(114), .d(8'h00));
tb.hm_put_byte(.addr(115), .d(8'h00));
tb.hm_put_byte(.addr(116), .d(8'h00));
tb.hm_put_byte(.addr(117), .d(8'h00));
tb.hm_put_byte(.addr(118), .d(8'h00));
tb.hm_put_byte(.addr(119), .d(8'h00));
tb.hm_put_byte(.addr(120), .d(8'h60));
tb.hm_put_byte(.addr(121), .d(8'hFF));
tb.hm_put_byte(.addr(122), .d(8'hFF));
tb.hm_put_byte(.addr(123), .d(8'hFF));
tb.hm_put_byte(.addr(124), .d(8'hFF));
tb.hm_put_byte(.addr(125), .d(8'hFF));
tb.hm_put_byte(.addr(126), .d(8'hFF));
tb.hm_put_byte(.addr(127), .d(8'hFF));
tb.hm_put_byte(.addr(128), .d(8'h0E));
tb.hm_put_byte(.addr(129), .d(8'h00));
tb.hm_put_byte(.addr(130), .d(8'h00));
tb.hm_put_byte(.addr(131), .d(8'h00));
tb.hm_put_byte(.addr(132), .d(8'h00));
tb.hm_put_byte(.addr(133), .d(8'h00));
tb.hm_put_byte(.addr(134), .d(8'h00));
tb.hm_put_byte(.addr(135), .d(8'h00));
tb.hm_put_byte(.addr(136), .d(8'h03));
tb.hm_put_byte(.addr(137), .d(8'h00));
tb.hm_put_byte(.addr(138), .d(8'h00));
tb.hm_put_byte(.addr(139), .d(8'h00));
tb.hm_put_byte(.addr(140), .d(8'h00));
tb.hm_put_byte(.addr(141), .d(8'h00));
tb.hm_put_byte(.addr(142), .d(8'h00));
tb.hm_put_byte(.addr(143), .d(8'h00));
tb.hm_put_byte(.addr(144), .d(8'h6F));
tb.hm_put_byte(.addr(145), .d(8'h00));
tb.hm_put_byte(.addr(146), .d(8'h00));
tb.hm_put_byte(.addr(147), .d(8'h00));
tb.hm_put_byte(.addr(148), .d(8'h00));
tb.hm_put_byte(.addr(149), .d(8'h00));
tb.hm_put_byte(.addr(150), .d(8'h00));
tb.hm_put_byte(.addr(151), .d(8'h00));
tb.hm_put_byte(.addr(152), .d(8'h79));
tb.hm_put_byte(.addr(153), .d(8'h00));
tb.hm_put_byte(.addr(154), .d(8'h00));
tb.hm_put_byte(.addr(155), .d(8'h00));
tb.hm_put_byte(.addr(156), .d(8'h00));
tb.hm_put_byte(.addr(157), .d(8'h00));
tb.hm_put_byte(.addr(158), .d(8'h00));
tb.hm_put_byte(.addr(159), .d(8'h00));
tb.hm_put_byte(.addr(160), .d(8'h83));
tb.hm_put_byte(.addr(161), .d(8'h00));
tb.hm_put_byte(.addr(162), .d(8'h00));
tb.hm_put_byte(.addr(163), .d(8'h00));
tb.hm_put_byte(.addr(164), .d(8'h00));
tb.hm_put_byte(.addr(165), .d(8'h00));
tb.hm_put_byte(.addr(166), .d(8'h00));
tb.hm_put_byte(.addr(167), .d(8'h00));
tb.hm_put_byte(.addr(168), .d(8'h8D));
tb.hm_put_byte(.addr(169), .d(8'h00));
tb.hm_put_byte(.addr(170), .d(8'h00));
tb.hm_put_byte(.addr(171), .d(8'h00));
tb.hm_put_byte(.addr(172), .d(8'h00));
tb.hm_put_byte(.addr(173), .d(8'h00));
tb.hm_put_byte(.addr(174), .d(8'h00));
tb.hm_put_byte(.addr(175), .d(8'h00));
tb.hm_put_byte(.addr(176), .d(8'h97));
tb.hm_put_byte(.addr(177), .d(8'h00));
tb.hm_put_byte(.addr(178), .d(8'h00));
tb.hm_put_byte(.addr(179), .d(8'h00));
tb.hm_put_byte(.addr(180), .d(8'h00));
tb.hm_put_byte(.addr(181), .d(8'h00));
tb.hm_put_byte(.addr(182), .d(8'h00));
tb.hm_put_byte(.addr(183), .d(8'h00));
tb.hm_put_byte(.addr(184), .d(8'h5F));
tb.hm_put_byte(.addr(185), .d(8'hFF));
tb.hm_put_byte(.addr(186), .d(8'hFF));
tb.hm_put_byte(.addr(187), .d(8'hFF));
tb.hm_put_byte(.addr(188), .d(8'hFF));
tb.hm_put_byte(.addr(189), .d(8'hFF));
tb.hm_put_byte(.addr(190), .d(8'hFF));
tb.hm_put_byte(.addr(191), .d(8'hFF));
tb.hm_put_byte(.addr(192), .d(8'h0D));
tb.hm_put_byte(.addr(193), .d(8'h00));
tb.hm_put_byte(.addr(194), .d(8'h00));
tb.hm_put_byte(.addr(195), .d(8'h00));
tb.hm_put_byte(.addr(196), .d(8'h00));
tb.hm_put_byte(.addr(197), .d(8'h00));
tb.hm_put_byte(.addr(198), .d(8'h00));
tb.hm_put_byte(.addr(199), .d(8'h00));
tb.hm_put_byte(.addr(200), .d(8'h00));
tb.hm_put_byte(.addr(201), .d(8'h00));
tb.hm_put_byte(.addr(202), .d(8'h00));
tb.hm_put_byte(.addr(203), .d(8'h00));
tb.hm_put_byte(.addr(204), .d(8'h00));
tb.hm_put_byte(.addr(205), .d(8'h00));
tb.hm_put_byte(.addr(206), .d(8'h00));
tb.hm_put_byte(.addr(207), .d(8'h00));
tb.hm_put_byte(.addr(208), .d(8'h70));
tb.hm_put_byte(.addr(209), .d(8'h00));
tb.hm_put_byte(.addr(210), .d(8'h00));
tb.hm_put_byte(.addr(211), .d(8'h00));
tb.hm_put_byte(.addr(212), .d(8'h00));
tb.hm_put_byte(.addr(213), .d(8'h00));
tb.hm_put_byte(.addr(214), .d(8'h00));
tb.hm_put_byte(.addr(215), .d(8'h00));
tb.hm_put_byte(.addr(216), .d(8'h7A));
tb.hm_put_byte(.addr(217), .d(8'h00));
tb.hm_put_byte(.addr(218), .d(8'h00));
tb.hm_put_byte(.addr(219), .d(8'h00));
tb.hm_put_byte(.addr(220), .d(8'h00));
tb.hm_put_byte(.addr(221), .d(8'h00));
tb.hm_put_byte(.addr(222), .d(8'h00));
tb.hm_put_byte(.addr(223), .d(8'h00));
tb.hm_put_byte(.addr(224), .d(8'h84));
tb.hm_put_byte(.addr(225), .d(8'h00));
tb.hm_put_byte(.addr(226), .d(8'h00));
tb.hm_put_byte(.addr(227), .d(8'h00));
tb.hm_put_byte(.addr(228), .d(8'h00));
tb.hm_put_byte(.addr(229), .d(8'h00));
tb.hm_put_byte(.addr(230), .d(8'h00));
tb.hm_put_byte(.addr(231), .d(8'h00));
tb.hm_put_byte(.addr(232), .d(8'h8E));
tb.hm_put_byte(.addr(233), .d(8'h00));
tb.hm_put_byte(.addr(234), .d(8'h00));
tb.hm_put_byte(.addr(235), .d(8'h00));
tb.hm_put_byte(.addr(236), .d(8'h00));
tb.hm_put_byte(.addr(237), .d(8'h00));
tb.hm_put_byte(.addr(238), .d(8'h00));
tb.hm_put_byte(.addr(239), .d(8'h00));
tb.hm_put_byte(.addr(240), .d(8'h98));
tb.hm_put_byte(.addr(241), .d(8'h00));
tb.hm_put_byte(.addr(242), .d(8'h00));
tb.hm_put_byte(.addr(243), .d(8'h00));
tb.hm_put_byte(.addr(244), .d(8'h00));
tb.hm_put_byte(.addr(245), .d(8'h00));
tb.hm_put_byte(.addr(246), .d(8'h00));
tb.hm_put_byte(.addr(247), .d(8'h00));
tb.hm_put_byte(.addr(248), .d(8'h5E));
tb.hm_put_byte(.addr(249), .d(8'hFF));
tb.hm_put_byte(.addr(250), .d(8'hFF));
tb.hm_put_byte(.addr(251), .d(8'hFF));
tb.hm_put_byte(.addr(252), .d(8'hFF));
tb.hm_put_byte(.addr(253), .d(8'hFF));
tb.hm_put_byte(.addr(254), .d(8'hFF));
tb.hm_put_byte(.addr(255), .d(8'hFF));
tb.hm_put_byte(.addr(256), .d(8'h2D));
tb.hm_put_byte(.addr(257), .d(8'h00));
tb.hm_put_byte(.addr(258), .d(8'h00));
tb.hm_put_byte(.addr(259), .d(8'h00));
tb.hm_put_byte(.addr(260), .d(8'h00));
tb.hm_put_byte(.addr(261), .d(8'h00));
tb.hm_put_byte(.addr(262), .d(8'h00));
tb.hm_put_byte(.addr(263), .d(8'h00));
tb.hm_put_byte(.addr(264), .d(8'h0C));
tb.hm_put_byte(.addr(265), .d(8'hFE));
tb.hm_put_byte(.addr(266), .d(8'hFF));
tb.hm_put_byte(.addr(267), .d(8'hFF));
tb.hm_put_byte(.addr(268), .d(8'hFF));
tb.hm_put_byte(.addr(269), .d(8'hFF));
tb.hm_put_byte(.addr(270), .d(8'hFF));
tb.hm_put_byte(.addr(271), .d(8'hFF));
tb.hm_put_byte(.addr(272), .d(8'hD2));
tb.hm_put_byte(.addr(273), .d(8'h00));
tb.hm_put_byte(.addr(274), .d(8'h00));
tb.hm_put_byte(.addr(275), .d(8'h00));
tb.hm_put_byte(.addr(276), .d(8'h00));
tb.hm_put_byte(.addr(277), .d(8'h00));
tb.hm_put_byte(.addr(278), .d(8'h00));
tb.hm_put_byte(.addr(279), .d(8'h00));
tb.hm_put_byte(.addr(280), .d(8'hDC));
tb.hm_put_byte(.addr(281), .d(8'h00));
tb.hm_put_byte(.addr(282), .d(8'h00));
tb.hm_put_byte(.addr(283), .d(8'h00));
tb.hm_put_byte(.addr(284), .d(8'h00));
tb.hm_put_byte(.addr(285), .d(8'h00));
tb.hm_put_byte(.addr(286), .d(8'h00));
tb.hm_put_byte(.addr(287), .d(8'h00));
tb.hm_put_byte(.addr(288), .d(8'hE6));
tb.hm_put_byte(.addr(289), .d(8'h00));
tb.hm_put_byte(.addr(290), .d(8'h00));
tb.hm_put_byte(.addr(291), .d(8'h00));
tb.hm_put_byte(.addr(292), .d(8'h00));
tb.hm_put_byte(.addr(293), .d(8'h00));
tb.hm_put_byte(.addr(294), .d(8'h00));
tb.hm_put_byte(.addr(295), .d(8'h00));
tb.hm_put_byte(.addr(296), .d(8'hF0));
tb.hm_put_byte(.addr(297), .d(8'h00));
tb.hm_put_byte(.addr(298), .d(8'h00));
tb.hm_put_byte(.addr(299), .d(8'h00));
tb.hm_put_byte(.addr(300), .d(8'h00));
tb.hm_put_byte(.addr(301), .d(8'h00));
tb.hm_put_byte(.addr(302), .d(8'h00));
tb.hm_put_byte(.addr(303), .d(8'h00));
tb.hm_put_byte(.addr(304), .d(8'hFA));
tb.hm_put_byte(.addr(305), .d(8'h00));
tb.hm_put_byte(.addr(306), .d(8'h00));
tb.hm_put_byte(.addr(307), .d(8'h00));
tb.hm_put_byte(.addr(308), .d(8'h00));
tb.hm_put_byte(.addr(309), .d(8'h00));
tb.hm_put_byte(.addr(310), .d(8'h00));
tb.hm_put_byte(.addr(311), .d(8'h00));
tb.hm_put_byte(.addr(312), .d(8'hFC));
tb.hm_put_byte(.addr(313), .d(8'hFE));
tb.hm_put_byte(.addr(314), .d(8'hFF));
tb.hm_put_byte(.addr(315), .d(8'hFF));
tb.hm_put_byte(.addr(316), .d(8'hFF));
tb.hm_put_byte(.addr(317), .d(8'hFF));
tb.hm_put_byte(.addr(318), .d(8'hFF));
tb.hm_put_byte(.addr(319), .d(8'hFF));
tb.hm_put_byte(.addr(320), .d(8'h33));
tb.hm_put_byte(.addr(321), .d(8'h00));
tb.hm_put_byte(.addr(322), .d(8'h00));
tb.hm_put_byte(.addr(323), .d(8'h00));
tb.hm_put_byte(.addr(324), .d(8'h00));
tb.hm_put_byte(.addr(325), .d(8'h00));
tb.hm_put_byte(.addr(326), .d(8'h00));
tb.hm_put_byte(.addr(327), .d(8'h00));
tb.hm_put_byte(.addr(328), .d(8'hF8));
tb.hm_put_byte(.addr(329), .d(8'hFD));
tb.hm_put_byte(.addr(330), .d(8'hFF));
tb.hm_put_byte(.addr(331), .d(8'hFF));
tb.hm_put_byte(.addr(332), .d(8'hFF));
tb.hm_put_byte(.addr(333), .d(8'hFF));
tb.hm_put_byte(.addr(334), .d(8'hFF));
tb.hm_put_byte(.addr(335), .d(8'hFF));
tb.hm_put_byte(.addr(336), .d(8'hD3));
tb.hm_put_byte(.addr(337), .d(8'h00));
tb.hm_put_byte(.addr(338), .d(8'h00));
tb.hm_put_byte(.addr(339), .d(8'h00));
tb.hm_put_byte(.addr(340), .d(8'h00));
tb.hm_put_byte(.addr(341), .d(8'h00));
tb.hm_put_byte(.addr(342), .d(8'h00));
tb.hm_put_byte(.addr(343), .d(8'h00));
tb.hm_put_byte(.addr(344), .d(8'hDD));
tb.hm_put_byte(.addr(345), .d(8'h00));
tb.hm_put_byte(.addr(346), .d(8'h00));
tb.hm_put_byte(.addr(347), .d(8'h00));
tb.hm_put_byte(.addr(348), .d(8'h00));
tb.hm_put_byte(.addr(349), .d(8'h00));
tb.hm_put_byte(.addr(350), .d(8'h00));
tb.hm_put_byte(.addr(351), .d(8'h00));
tb.hm_put_byte(.addr(352), .d(8'hE7));
tb.hm_put_byte(.addr(353), .d(8'h00));
tb.hm_put_byte(.addr(354), .d(8'h00));
tb.hm_put_byte(.addr(355), .d(8'h00));
tb.hm_put_byte(.addr(356), .d(8'h00));
tb.hm_put_byte(.addr(357), .d(8'h00));
tb.hm_put_byte(.addr(358), .d(8'h00));
tb.hm_put_byte(.addr(359), .d(8'h00));
tb.hm_put_byte(.addr(360), .d(8'hF1));
tb.hm_put_byte(.addr(361), .d(8'h00));
tb.hm_put_byte(.addr(362), .d(8'h00));
tb.hm_put_byte(.addr(363), .d(8'h00));
tb.hm_put_byte(.addr(364), .d(8'h00));
tb.hm_put_byte(.addr(365), .d(8'h00));
tb.hm_put_byte(.addr(366), .d(8'h00));
tb.hm_put_byte(.addr(367), .d(8'h00));
tb.hm_put_byte(.addr(368), .d(8'h97));
tb.hm_put_byte(.addr(369), .d(8'h00));
tb.hm_put_byte(.addr(370), .d(8'h00));
tb.hm_put_byte(.addr(371), .d(8'h00));
tb.hm_put_byte(.addr(372), .d(8'h00));
tb.hm_put_byte(.addr(373), .d(8'h00));
tb.hm_put_byte(.addr(374), .d(8'h00));
tb.hm_put_byte(.addr(375), .d(8'h00));
tb.hm_put_byte(.addr(376), .d(8'hFB));
tb.hm_put_byte(.addr(377), .d(8'hFE));
tb.hm_put_byte(.addr(378), .d(8'hFF));
tb.hm_put_byte(.addr(379), .d(8'hFF));
tb.hm_put_byte(.addr(380), .d(8'hFF));
tb.hm_put_byte(.addr(381), .d(8'hFF));
tb.hm_put_byte(.addr(382), .d(8'hFF));
tb.hm_put_byte(.addr(383), .d(8'hFF));
