-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.UtilStr_pkg.all;
use work.UtilConv_pkg.all;

entity Profiler is
  generic (
    PROBE_COUNT_WIDTH : positive;
    OUT_COUNT_WIDTH   : positive
  );
  port (
    pcd_clk         : in  std_logic;
    pcd_reset       : in  std_logic;
    probe_valid     : in  std_logic;
    probe_ready     : in  std_logic;
    probe_last      : in  std_logic;
    probe_count     : in  std_logic_vector(PROBE_COUNT_WIDTH-1 downto 0) := std_logic_vector(to_unsigned(1, PROBE_COUNT_WIDTH));
    enable          : in  std_logic;
    clear           : in  std_logic;
    count_elements  : out std_logic_vector(OUT_COUNT_WIDTH-1 downto 0);
    count_valids    : out std_logic_vector(OUT_COUNT_WIDTH-1 downto 0);
    count_readies   : out std_logic_vector(OUT_COUNT_WIDTH-1 downto 0);
    count_transfers : out std_logic_vector(OUT_COUNT_WIDTH-1 downto 0);
    count_packets   : out std_logic_vector(OUT_COUNT_WIDTH-1 downto 0);
    count_cycles    : out std_logic_vector(OUT_COUNT_WIDTH-1 downto 0)
  );
end Profiler;

architecture Behavioral of Profiler is
begin

process(pcd_clk) is
  constant ZERO_COUNT : unsigned(OUT_COUNT_WIDTH-1 downto 0) := to_unsigned(0, OUT_COUNT_WIDTH);
  variable elements   : unsigned(OUT_COUNT_WIDTH-1 downto 0) := ZERO_COUNT;
  variable valids     : unsigned(OUT_COUNT_WIDTH-1 downto 0) := ZERO_COUNT;
  variable readies    : unsigned(OUT_COUNT_WIDTH-1 downto 0) := ZERO_COUNT;
  variable transfers  : unsigned(OUT_COUNT_WIDTH-1 downto 0) := ZERO_COUNT;
  variable packets    : unsigned(OUT_COUNT_WIDTH-1 downto 0) := ZERO_COUNT;
  variable cycles     : unsigned(OUT_COUNT_WIDTH-1 downto 0) := ZERO_COUNT;
begin
  if rising_edge(pcd_clk) then
    if (enable = '1') then
      if (probe_valid = '1') then
        valids := valids + 1;
      end if;
      if (probe_ready = '1') then
        readies := readies + 1;
      end if;
      if (probe_valid = '1') and (probe_ready = '1') then
        transfers := transfers + 1;
      end if;
      if (probe_valid = '1') and (probe_ready = '1') and (probe_last = '1') then
        packets := packets + 1;
      end if;

      cycles := cycles + 1;
    end if;

    if (pcd_reset = '1') or (clear = '1') then
      elements  := ZERO_COUNT;
      valids    := ZERO_COUNT;
      readies   := ZERO_COUNT;
      transfers := ZERO_COUNT;
      packets   := ZERO_COUNT;
      cycles    := ZERO_COUNT;
    end if;

    count_elements  <= std_logic_vector(elements);
    count_valids    <= std_logic_vector(valids);
    count_readies   <= std_logic_vector(readies);
    count_transfers <= std_logic_vector(transfers);
    count_packets   <= std_logic_vector(packets);
    count_cycles    <= std_logic_vector(cycles);
  end if;

end process;

end architecture;
