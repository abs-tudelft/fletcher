tb.hm_put_byte(.addr(0), .d(8'h00));
tb.hm_put_byte(.addr(1), .d(8'h00));
tb.hm_put_byte(.addr(2), .d(8'h00));
tb.hm_put_byte(.addr(3), .d(8'h00));
tb.hm_put_byte(.addr(4), .d(8'h02));
tb.hm_put_byte(.addr(5), .d(8'h00));
tb.hm_put_byte(.addr(6), .d(8'h00));
tb.hm_put_byte(.addr(7), .d(8'h00));
tb.hm_put_byte(.addr(8), .d(8'h04));
tb.hm_put_byte(.addr(9), .d(8'h00));
tb.hm_put_byte(.addr(10), .d(8'h00));
tb.hm_put_byte(.addr(11), .d(8'h00));
tb.hm_put_byte(.addr(12), .d(8'h06));
tb.hm_put_byte(.addr(13), .d(8'h00));
tb.hm_put_byte(.addr(14), .d(8'h00));
tb.hm_put_byte(.addr(15), .d(8'h00));
tb.hm_put_byte(.addr(16), .d(8'h08));
tb.hm_put_byte(.addr(17), .d(8'h00));
tb.hm_put_byte(.addr(18), .d(8'h00));
tb.hm_put_byte(.addr(19), .d(8'h00));
tb.hm_put_byte(.addr(20), .d(8'h0A));
tb.hm_put_byte(.addr(21), .d(8'h00));
tb.hm_put_byte(.addr(22), .d(8'h00));
tb.hm_put_byte(.addr(23), .d(8'h00));
tb.hm_put_byte(.addr(24), .d(8'h00));
tb.hm_put_byte(.addr(25), .d(8'h00));
tb.hm_put_byte(.addr(26), .d(8'h00));
tb.hm_put_byte(.addr(27), .d(8'h00));
tb.hm_put_byte(.addr(28), .d(8'h00));
tb.hm_put_byte(.addr(29), .d(8'h00));
tb.hm_put_byte(.addr(30), .d(8'h00));
tb.hm_put_byte(.addr(31), .d(8'h00));
tb.hm_put_byte(.addr(32), .d(8'h00));
tb.hm_put_byte(.addr(33), .d(8'h00));
tb.hm_put_byte(.addr(34), .d(8'h00));
tb.hm_put_byte(.addr(35), .d(8'h00));
tb.hm_put_byte(.addr(36), .d(8'h00));
tb.hm_put_byte(.addr(37), .d(8'h00));
tb.hm_put_byte(.addr(38), .d(8'h00));
tb.hm_put_byte(.addr(39), .d(8'h00));
tb.hm_put_byte(.addr(40), .d(8'h00));
tb.hm_put_byte(.addr(41), .d(8'h00));
tb.hm_put_byte(.addr(42), .d(8'h00));
tb.hm_put_byte(.addr(43), .d(8'h00));
tb.hm_put_byte(.addr(44), .d(8'h00));
tb.hm_put_byte(.addr(45), .d(8'h00));
tb.hm_put_byte(.addr(46), .d(8'h00));
tb.hm_put_byte(.addr(47), .d(8'h00));
tb.hm_put_byte(.addr(48), .d(8'h00));
tb.hm_put_byte(.addr(49), .d(8'h00));
tb.hm_put_byte(.addr(50), .d(8'h00));
tb.hm_put_byte(.addr(51), .d(8'h00));
tb.hm_put_byte(.addr(52), .d(8'h00));
tb.hm_put_byte(.addr(53), .d(8'h00));
tb.hm_put_byte(.addr(54), .d(8'h00));
tb.hm_put_byte(.addr(55), .d(8'h00));
tb.hm_put_byte(.addr(56), .d(8'h00));
tb.hm_put_byte(.addr(57), .d(8'h00));
tb.hm_put_byte(.addr(58), .d(8'h00));
tb.hm_put_byte(.addr(59), .d(8'h00));
tb.hm_put_byte(.addr(60), .d(8'h00));
tb.hm_put_byte(.addr(61), .d(8'h00));
tb.hm_put_byte(.addr(62), .d(8'h00));
tb.hm_put_byte(.addr(63), .d(8'h00));
tb.hm_put_byte(.addr(64), .d(8'h0C));
tb.hm_put_byte(.addr(65), .d(8'h00));
tb.hm_put_byte(.addr(66), .d(8'h00));
tb.hm_put_byte(.addr(67), .d(8'h00));
tb.hm_put_byte(.addr(68), .d(8'h00));
tb.hm_put_byte(.addr(69), .d(8'h00));
tb.hm_put_byte(.addr(70), .d(8'h00));
tb.hm_put_byte(.addr(71), .d(8'h00));
tb.hm_put_byte(.addr(72), .d(8'h06));
tb.hm_put_byte(.addr(73), .d(8'h00));
tb.hm_put_byte(.addr(74), .d(8'h00));
tb.hm_put_byte(.addr(75), .d(8'h00));
tb.hm_put_byte(.addr(76), .d(8'h00));
tb.hm_put_byte(.addr(77), .d(8'h00));
tb.hm_put_byte(.addr(78), .d(8'h00));
tb.hm_put_byte(.addr(79), .d(8'h00));
tb.hm_put_byte(.addr(80), .d(8'h0E));
tb.hm_put_byte(.addr(81), .d(8'h00));
tb.hm_put_byte(.addr(82), .d(8'h00));
tb.hm_put_byte(.addr(83), .d(8'h00));
tb.hm_put_byte(.addr(84), .d(8'h00));
tb.hm_put_byte(.addr(85), .d(8'h00));
tb.hm_put_byte(.addr(86), .d(8'h00));
tb.hm_put_byte(.addr(87), .d(8'h00));
tb.hm_put_byte(.addr(88), .d(8'h03));
tb.hm_put_byte(.addr(89), .d(8'h00));
tb.hm_put_byte(.addr(90), .d(8'h00));
tb.hm_put_byte(.addr(91), .d(8'h00));
tb.hm_put_byte(.addr(92), .d(8'h00));
tb.hm_put_byte(.addr(93), .d(8'h00));
tb.hm_put_byte(.addr(94), .d(8'h00));
tb.hm_put_byte(.addr(95), .d(8'h00));
tb.hm_put_byte(.addr(96), .d(8'h0D));
tb.hm_put_byte(.addr(97), .d(8'h00));
tb.hm_put_byte(.addr(98), .d(8'h00));
tb.hm_put_byte(.addr(99), .d(8'h00));
tb.hm_put_byte(.addr(100), .d(8'h00));
tb.hm_put_byte(.addr(101), .d(8'h00));
tb.hm_put_byte(.addr(102), .d(8'h00));
tb.hm_put_byte(.addr(103), .d(8'h00));
tb.hm_put_byte(.addr(104), .d(8'h00));
tb.hm_put_byte(.addr(105), .d(8'h00));
tb.hm_put_byte(.addr(106), .d(8'h00));
tb.hm_put_byte(.addr(107), .d(8'h00));
tb.hm_put_byte(.addr(108), .d(8'h00));
tb.hm_put_byte(.addr(109), .d(8'h00));
tb.hm_put_byte(.addr(110), .d(8'h00));
tb.hm_put_byte(.addr(111), .d(8'h00));
tb.hm_put_byte(.addr(112), .d(8'h2D));
tb.hm_put_byte(.addr(113), .d(8'h00));
tb.hm_put_byte(.addr(114), .d(8'h00));
tb.hm_put_byte(.addr(115), .d(8'h00));
tb.hm_put_byte(.addr(116), .d(8'h00));
tb.hm_put_byte(.addr(117), .d(8'h00));
tb.hm_put_byte(.addr(118), .d(8'h00));
tb.hm_put_byte(.addr(119), .d(8'h00));
tb.hm_put_byte(.addr(120), .d(8'h0C));
tb.hm_put_byte(.addr(121), .d(8'hFE));
tb.hm_put_byte(.addr(122), .d(8'hFF));
tb.hm_put_byte(.addr(123), .d(8'hFF));
tb.hm_put_byte(.addr(124), .d(8'hFF));
tb.hm_put_byte(.addr(125), .d(8'hFF));
tb.hm_put_byte(.addr(126), .d(8'hFF));
tb.hm_put_byte(.addr(127), .d(8'hFF));
tb.hm_put_byte(.addr(128), .d(8'h33));
tb.hm_put_byte(.addr(129), .d(8'h00));
tb.hm_put_byte(.addr(130), .d(8'h00));
tb.hm_put_byte(.addr(131), .d(8'h00));
tb.hm_put_byte(.addr(132), .d(8'h00));
tb.hm_put_byte(.addr(133), .d(8'h00));
tb.hm_put_byte(.addr(134), .d(8'h00));
tb.hm_put_byte(.addr(135), .d(8'h00));
tb.hm_put_byte(.addr(136), .d(8'hF8));
tb.hm_put_byte(.addr(137), .d(8'hFD));
tb.hm_put_byte(.addr(138), .d(8'hFF));
tb.hm_put_byte(.addr(139), .d(8'hFF));
tb.hm_put_byte(.addr(140), .d(8'hFF));
tb.hm_put_byte(.addr(141), .d(8'hFF));
tb.hm_put_byte(.addr(142), .d(8'hFF));
tb.hm_put_byte(.addr(143), .d(8'hFF));
tb.hm_put_byte(.addr(144), .d(8'h00));
tb.hm_put_byte(.addr(145), .d(8'h00));
tb.hm_put_byte(.addr(146), .d(8'h00));
tb.hm_put_byte(.addr(147), .d(8'h00));
tb.hm_put_byte(.addr(148), .d(8'h00));
tb.hm_put_byte(.addr(149), .d(8'h00));
tb.hm_put_byte(.addr(150), .d(8'h00));
tb.hm_put_byte(.addr(151), .d(8'h00));
tb.hm_put_byte(.addr(152), .d(8'h00));
tb.hm_put_byte(.addr(153), .d(8'h00));
tb.hm_put_byte(.addr(154), .d(8'h00));
tb.hm_put_byte(.addr(155), .d(8'h00));
tb.hm_put_byte(.addr(156), .d(8'h00));
tb.hm_put_byte(.addr(157), .d(8'h00));
tb.hm_put_byte(.addr(158), .d(8'h00));
tb.hm_put_byte(.addr(159), .d(8'h00));
tb.hm_put_byte(.addr(160), .d(8'h00));
tb.hm_put_byte(.addr(161), .d(8'h00));
tb.hm_put_byte(.addr(162), .d(8'h00));
tb.hm_put_byte(.addr(163), .d(8'h00));
tb.hm_put_byte(.addr(164), .d(8'h00));
tb.hm_put_byte(.addr(165), .d(8'h00));
tb.hm_put_byte(.addr(166), .d(8'h00));
tb.hm_put_byte(.addr(167), .d(8'h00));
tb.hm_put_byte(.addr(168), .d(8'h00));
tb.hm_put_byte(.addr(169), .d(8'h00));
tb.hm_put_byte(.addr(170), .d(8'h00));
tb.hm_put_byte(.addr(171), .d(8'h00));
tb.hm_put_byte(.addr(172), .d(8'h00));
tb.hm_put_byte(.addr(173), .d(8'h00));
tb.hm_put_byte(.addr(174), .d(8'h00));
tb.hm_put_byte(.addr(175), .d(8'h00));
tb.hm_put_byte(.addr(176), .d(8'h00));
tb.hm_put_byte(.addr(177), .d(8'h00));
tb.hm_put_byte(.addr(178), .d(8'h00));
tb.hm_put_byte(.addr(179), .d(8'h00));
tb.hm_put_byte(.addr(180), .d(8'h00));
tb.hm_put_byte(.addr(181), .d(8'h00));
tb.hm_put_byte(.addr(182), .d(8'h00));
tb.hm_put_byte(.addr(183), .d(8'h00));
tb.hm_put_byte(.addr(184), .d(8'h00));
tb.hm_put_byte(.addr(185), .d(8'h00));
tb.hm_put_byte(.addr(186), .d(8'h00));
tb.hm_put_byte(.addr(187), .d(8'h00));
tb.hm_put_byte(.addr(188), .d(8'h00));
tb.hm_put_byte(.addr(189), .d(8'h00));
tb.hm_put_byte(.addr(190), .d(8'h00));
tb.hm_put_byte(.addr(191), .d(8'h00));
