tb.hm_put_byte(.addr(0), .d(8'h00));
tb.hm_put_byte(.addr(1), .d(8'h00));
tb.hm_put_byte(.addr(2), .d(8'h00));
tb.hm_put_byte(.addr(3), .d(8'h00));
tb.hm_put_byte(.addr(4), .d(8'h02));
tb.hm_put_byte(.addr(5), .d(8'h00));
tb.hm_put_byte(.addr(6), .d(8'h00));
tb.hm_put_byte(.addr(7), .d(8'h00));
tb.hm_put_byte(.addr(8), .d(8'h04));
tb.hm_put_byte(.addr(9), .d(8'h00));
tb.hm_put_byte(.addr(10), .d(8'h00));
tb.hm_put_byte(.addr(11), .d(8'h00));
tb.hm_put_byte(.addr(12), .d(8'h06));
tb.hm_put_byte(.addr(13), .d(8'h00));
tb.hm_put_byte(.addr(14), .d(8'h00));
tb.hm_put_byte(.addr(15), .d(8'h00));
tb.hm_put_byte(.addr(16), .d(8'h08));
tb.hm_put_byte(.addr(17), .d(8'h00));
tb.hm_put_byte(.addr(18), .d(8'h00));
tb.hm_put_byte(.addr(19), .d(8'h00));
tb.hm_put_byte(.addr(20), .d(8'h00));
tb.hm_put_byte(.addr(21), .d(8'h00));
tb.hm_put_byte(.addr(22), .d(8'h00));
tb.hm_put_byte(.addr(23), .d(8'h00));
tb.hm_put_byte(.addr(24), .d(8'h00));
tb.hm_put_byte(.addr(25), .d(8'h00));
tb.hm_put_byte(.addr(26), .d(8'h00));
tb.hm_put_byte(.addr(27), .d(8'h00));
tb.hm_put_byte(.addr(28), .d(8'h00));
tb.hm_put_byte(.addr(29), .d(8'h00));
tb.hm_put_byte(.addr(30), .d(8'h00));
tb.hm_put_byte(.addr(31), .d(8'h00));
tb.hm_put_byte(.addr(32), .d(8'h00));
tb.hm_put_byte(.addr(33), .d(8'h00));
tb.hm_put_byte(.addr(34), .d(8'h00));
tb.hm_put_byte(.addr(35), .d(8'h00));
tb.hm_put_byte(.addr(36), .d(8'h00));
tb.hm_put_byte(.addr(37), .d(8'h00));
tb.hm_put_byte(.addr(38), .d(8'h00));
tb.hm_put_byte(.addr(39), .d(8'h00));
tb.hm_put_byte(.addr(40), .d(8'h00));
tb.hm_put_byte(.addr(41), .d(8'h00));
tb.hm_put_byte(.addr(42), .d(8'h00));
tb.hm_put_byte(.addr(43), .d(8'h00));
tb.hm_put_byte(.addr(44), .d(8'h00));
tb.hm_put_byte(.addr(45), .d(8'h00));
tb.hm_put_byte(.addr(46), .d(8'h00));
tb.hm_put_byte(.addr(47), .d(8'h00));
tb.hm_put_byte(.addr(48), .d(8'h00));
tb.hm_put_byte(.addr(49), .d(8'h00));
tb.hm_put_byte(.addr(50), .d(8'h00));
tb.hm_put_byte(.addr(51), .d(8'h00));
tb.hm_put_byte(.addr(52), .d(8'h00));
tb.hm_put_byte(.addr(53), .d(8'h00));
tb.hm_put_byte(.addr(54), .d(8'h00));
tb.hm_put_byte(.addr(55), .d(8'h00));
tb.hm_put_byte(.addr(56), .d(8'h00));
tb.hm_put_byte(.addr(57), .d(8'h00));
tb.hm_put_byte(.addr(58), .d(8'h00));
tb.hm_put_byte(.addr(59), .d(8'h00));
tb.hm_put_byte(.addr(60), .d(8'h00));
tb.hm_put_byte(.addr(61), .d(8'h00));
tb.hm_put_byte(.addr(62), .d(8'h00));
tb.hm_put_byte(.addr(63), .d(8'h00));
tb.hm_put_byte(.addr(64), .d(8'h33));
tb.hm_put_byte(.addr(65), .d(8'h33));
tb.hm_put_byte(.addr(66), .d(8'h33));
tb.hm_put_byte(.addr(67), .d(8'h33));
tb.hm_put_byte(.addr(68), .d(8'h33));
tb.hm_put_byte(.addr(69), .d(8'h33));
tb.hm_put_byte(.addr(70), .d(8'hF3));
tb.hm_put_byte(.addr(71), .d(8'h3F));
tb.hm_put_byte(.addr(72), .d(8'h33));
tb.hm_put_byte(.addr(73), .d(8'h33));
tb.hm_put_byte(.addr(74), .d(8'h33));
tb.hm_put_byte(.addr(75), .d(8'h33));
tb.hm_put_byte(.addr(76), .d(8'h33));
tb.hm_put_byte(.addr(77), .d(8'h33));
tb.hm_put_byte(.addr(78), .d(8'hE3));
tb.hm_put_byte(.addr(79), .d(8'h3F));
tb.hm_put_byte(.addr(80), .d(8'h66));
tb.hm_put_byte(.addr(81), .d(8'h66));
tb.hm_put_byte(.addr(82), .d(8'h66));
tb.hm_put_byte(.addr(83), .d(8'h66));
tb.hm_put_byte(.addr(84), .d(8'h66));
tb.hm_put_byte(.addr(85), .d(8'h66));
tb.hm_put_byte(.addr(86), .d(8'hF6));
tb.hm_put_byte(.addr(87), .d(8'h3F));
tb.hm_put_byte(.addr(88), .d(8'h33));
tb.hm_put_byte(.addr(89), .d(8'h33));
tb.hm_put_byte(.addr(90), .d(8'h33));
tb.hm_put_byte(.addr(91), .d(8'h33));
tb.hm_put_byte(.addr(92), .d(8'h33));
tb.hm_put_byte(.addr(93), .d(8'h33));
tb.hm_put_byte(.addr(94), .d(8'hD3));
tb.hm_put_byte(.addr(95), .d(8'h3F));
tb.hm_put_byte(.addr(96), .d(8'h00));
tb.hm_put_byte(.addr(97), .d(8'h00));
tb.hm_put_byte(.addr(98), .d(8'h00));
tb.hm_put_byte(.addr(99), .d(8'h00));
tb.hm_put_byte(.addr(100), .d(8'h00));
tb.hm_put_byte(.addr(101), .d(8'h00));
tb.hm_put_byte(.addr(102), .d(8'h12));
tb.hm_put_byte(.addr(103), .d(8'h40));
tb.hm_put_byte(.addr(104), .d(8'h33));
tb.hm_put_byte(.addr(105), .d(8'h33));
tb.hm_put_byte(.addr(106), .d(8'h33));
tb.hm_put_byte(.addr(107), .d(8'h33));
tb.hm_put_byte(.addr(108), .d(8'h33));
tb.hm_put_byte(.addr(109), .d(8'h33));
tb.hm_put_byte(.addr(110), .d(8'hF3));
tb.hm_put_byte(.addr(111), .d(8'hBF));
tb.hm_put_byte(.addr(112), .d(8'h66));
tb.hm_put_byte(.addr(113), .d(8'h66));
tb.hm_put_byte(.addr(114), .d(8'h66));
tb.hm_put_byte(.addr(115), .d(8'h66));
tb.hm_put_byte(.addr(116), .d(8'h66));
tb.hm_put_byte(.addr(117), .d(8'h66));
tb.hm_put_byte(.addr(118), .d(8'h14));
tb.hm_put_byte(.addr(119), .d(8'h40));
tb.hm_put_byte(.addr(120), .d(8'hCD));
tb.hm_put_byte(.addr(121), .d(8'hCC));
tb.hm_put_byte(.addr(122), .d(8'hCC));
tb.hm_put_byte(.addr(123), .d(8'hCC));
tb.hm_put_byte(.addr(124), .d(8'hCC));
tb.hm_put_byte(.addr(125), .d(8'hCC));
tb.hm_put_byte(.addr(126), .d(8'hF4));
tb.hm_put_byte(.addr(127), .d(8'hBF));
