-- Copyright 2018 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.

-- This file was automatically generated by FletchGen. Modify this file
-- at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;

library work;
use work.Arrow.all;
use work.Columns.all;
use work.Interconnect.all;
use work.Wrapper.all;

entity stringwrite_wrapper is
  generic(
    BUS_ADDR_WIDTH                             : natural;
    BUS_DATA_WIDTH                             : natural;
    BUS_STROBE_WIDTH                           : natural;
    BUS_LEN_WIDTH                              : natural;
    BUS_BURST_STEP_LEN                         : natural;
    BUS_BURST_MAX_LEN                          : natural;
    ---------------------------------------------------------------------------
    INDEX_WIDTH                                : natural;
    ---------------------------------------------------------------------------
    NUM_ARROW_BUFFERS                          : natural;
    NUM_REGS                                   : natural;
    NUM_USER_REGS                              : natural;
    REG_WIDTH                                  : natural;
    ---------------------------------------------------------------------------
    TAG_WIDTH                                  : natural
  );
  port(
    acc_reset                                  : in std_logic;
    bus_clk                                    : in std_logic;
    bus_reset                                  : in std_logic;
    acc_clk                                    : in std_logic;
    ---------------------------------------------------------------------------
    mst_rreq_valid                             : out std_logic;
    mst_rreq_ready                             : in std_logic;
    mst_rreq_addr                              : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    mst_rreq_len                               : out std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
    ---------------------------------------------------------------------------
    mst_rdat_valid                             : in std_logic;
    mst_rdat_ready                             : out std_logic;
    mst_rdat_data                              : in std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
    mst_rdat_last                              : in std_logic;
    ---------------------------------------------------------------------------
    mst_wreq_valid                             : out std_logic;
    mst_wreq_len                               : out std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
    mst_wreq_addr                              : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    mst_wreq_ready                             : in std_logic;
    ---------------------------------------------------------------------------
    mst_wdat_valid                             : out std_logic;
    mst_wdat_ready                             : in std_logic;
    mst_wdat_data                              : out std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
    mst_wdat_strobe                            : out std_logic_vector(BUS_STROBE_WIDTH-1 downto 0);
    mst_wdat_last                              : out std_logic;
    ---------------------------------------------------------------------------
    regs_in                                    : in std_logic_vector(NUM_REGS*REG_WIDTH-1 downto 0);
    regs_out                                   : out std_logic_vector(NUM_REGS*REG_WIDTH-1 downto 0);
    regs_out_en                                : out std_logic_vector(NUM_REGS-1 downto 0)
  );
end stringwrite_wrapper;

architecture Implementation of stringwrite_wrapper is

  -----------------------------------------------------------------------------
  -- Hardware Accelerated Function component.
  -- This component should be implemented by the user.
  component stringwrite_usercore is
    generic(
      NUM_USER_REGS                              : natural;
      TAG_WIDTH                                  : natural;
      BUS_ADDR_WIDTH                             : natural;
      INDEX_WIDTH                                : natural;
      REG_WIDTH                                  : natural
    );
    port(
      -------------------------------------------------------------------------
      acc_reset                                  : in std_logic;
      acc_clk                                    : in std_logic;
      -------------------------------------------------------------------------
      Str_in_values_in_count                     : out std_logic_vector(6 downto 0);
      Str_in_values_in_data                      : out std_logic_vector(511 downto 0);
      Str_in_values_in_dvalid                    : out std_logic;
      Str_in_values_in_last                      : out std_logic;
      Str_in_values_in_valid                     : out std_logic;
      Str_in_values_in_ready                     : in std_logic;
      -------------------------------------------------------------------------
      Str_in_length                              : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      Str_in_last                                : out std_logic;
      Str_in_valid                               : out std_logic;
      Str_in_dvalid                              : out std_logic;
      Str_in_ready                               : in std_logic;
      -------------------------------------------------------------------------
      Str_cmd_firstIdx                           : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      Str_cmd_lastIdx                            : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      Str_cmd_tag                                : out std_logic_vector(TAG_WIDTH-1 downto 0);
      Str_cmd_Str_offsets_addr                   : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      Str_cmd_Str_values_addr                    : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      Str_cmd_valid                              : out std_logic;
      Str_cmd_ready                              : in std_logic;
      -------------------------------------------------------------------------
      Str_unl_valid                              : in std_logic;
      Str_unl_ready                              : out std_logic;
      Str_unl_tag                                : in std_logic_vector(TAG_WIDTH-1 downto 0);
      -------------------------------------------------------------------------
      ctrl_done                                  : out std_logic;
      ctrl_busy                                  : out std_logic;
      ctrl_idle                                  : out std_logic;
      ctrl_reset                                 : in std_logic;
      ctrl_stop                                  : in std_logic;
      ctrl_start                                 : in std_logic;
      -------------------------------------------------------------------------
      reg_Str_offsets_addr                       : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      reg_Str_values_addr                        : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      -------------------------------------------------------------------------
      idx_first                                  : in std_logic_vector(REG_WIDTH-1 downto 0);
      idx_last                                   : in std_logic_vector(REG_WIDTH-1 downto 0);
      reg_return0                                : out std_logic_vector(REG_WIDTH-1 downto 0);
      reg_return1                                : out std_logic_vector(REG_WIDTH-1 downto 0);
      -------------------------------------------------------------------------
      regs_in                                    : in std_logic_vector(NUM_USER_REGS*REG_WIDTH-1 downto 0);
      regs_out                                   : out std_logic_vector(NUM_USER_REGS*REG_WIDTH-1 downto 0);
      regs_out_en                                : out std_logic_vector(NUM_USER_REGS-1 downto 0)
    );
  end component;
  -----------------------------------------------------------------------------
  signal uctrl_done                            : std_logic;
  signal uctrl_busy                            : std_logic;
  signal uctrl_idle                            : std_logic;
  signal uctrl_reset                           : std_logic;
  signal uctrl_stop                            : std_logic;
  signal uctrl_start                           : std_logic;
  signal uctrl_control                         : std_logic_vector(REG_WIDTH-1 downto 0);
  signal uctrl_status                          : std_logic_vector(REG_WIDTH-1 downto 0);
  -----------------------------------------------------------------------------
  signal s_Str_bus_wdat_last                   : std_logic;
  signal s_Str_bus_wdat_strobe                 : std_logic_vector(BUS_STROBE_WIDTH-1 downto 0);
  signal s_Str_bus_wdat_data                   : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal s_Str_bus_wdat_ready                  : std_logic;
  signal s_Str_bus_wdat_valid                  : std_logic;
  signal s_Str_bus_wreq_addr                   : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_Str_bus_wreq_len                    : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal s_Str_bus_wreq_ready                  : std_logic;
  signal s_Str_bus_wreq_valid                  : std_logic;
  -----------------------------------------------------------------------------
  signal s_Str_cmd_valid                       : std_logic;
  signal s_Str_cmd_ready                       : std_logic;
  signal s_Str_cmd_firstIdx                    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_Str_cmd_lastIdx                     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_Str_cmd_ctrl                        : std_logic_vector(2*BUS_ADDR_WIDTH-1 downto 0);
  signal s_Str_cmd_tag                         : std_logic_vector(TAG_WIDTH-1 downto 0);
  -----------------------------------------------------------------------------
  signal s_Str_in_valid                        : std_logic_vector(1 downto 0);
  signal s_Str_in_ready                        : std_logic_vector(1 downto 0);
  signal s_Str_in_last                         : std_logic_vector(1 downto 0);
  signal s_Str_in_dvalid                       : std_logic_vector(1 downto 0);
  signal s_Str_in_data                         : std_logic_vector(INDEX_WIDTH+518 downto 0);
  -----------------------------------------------------------------------------
  signal s_Str_unl_valid                       : std_logic;
  signal s_Str_unl_ready                       : std_logic;
  signal s_Str_unl_tag                         : std_logic_vector(TAG_WIDTH-1 downto 0);
  -----------------------------------------------------------------------------
  signal s_bsv_wreq_len                        : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal s_bsv_wreq_valid                      : std_logic_vector(0 downto 0);
  signal s_bsv_wreq_ready                      : std_logic_vector(0 downto 0);
  signal s_bsv_wreq_addr                       : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  -----------------------------------------------------------------------------
  signal s_bsv_wdat_valid                      : std_logic_vector(0 downto 0);
  signal s_bsv_wdat_last                       : std_logic_vector(0 downto 0);
  signal s_bsv_wdat_strobe                     : std_logic_vector(BUS_STROBE_WIDTH-1 downto 0);
  signal s_bsv_wdat_data                       : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal s_bsv_wdat_ready                      : std_logic_vector(0 downto 0);
  -----------------------------------------------------------------------------
  signal s_regs_out_en                         : std_logic_vector(NUM_USER_REGS-1 downto 0);
  signal s_regs_out                            : std_logic_vector(NUM_USER_REGS*REG_WIDTH-1 downto 0);
  signal s_regs_in                             : std_logic_vector(NUM_USER_REGS*REG_WIDTH-1 downto 0);

begin
  -- ColumnWriter instance generated from Arrow schema field:
  -- Str: string not null
  Str_write_inst: ColumnWriter
    generic map (
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH                            => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH                           => BUS_DATA_WIDTH,
      BUS_STROBE_WIDTH                         => BUS_STROBE_WIDTH,
      BUS_BURST_STEP_LEN                       => BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN                        => BUS_BURST_MAX_LEN,
      INDEX_WIDTH                              => INDEX_WIDTH,
      CFG                                      => "listprim(8;epc=64)",
      CMD_TAG_ENABLE                           => true,
      CMD_TAG_WIDTH                            => TAG_WIDTH
    )
    port map (
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      cmd_valid                                => s_Str_cmd_valid,
      cmd_ready                                => s_Str_cmd_ready,
      cmd_firstIdx                             => s_Str_cmd_firstIdx,
      cmd_lastIdx                              => s_Str_cmd_lastIdx,
      cmd_ctrl                                 => s_Str_cmd_ctrl,
      cmd_tag                                  => s_Str_cmd_tag,
      in_valid                                 => s_Str_in_valid,
      in_ready                                 => s_Str_in_ready,
      in_last                                  => s_Str_in_last,
      in_data                                  => s_Str_in_data,
      in_dvalid                                => s_Str_in_dvalid,
      bus_wreq_valid                           => s_Str_bus_wreq_valid,
      bus_wreq_ready                           => s_Str_bus_wreq_ready,
      bus_wreq_addr                            => s_Str_bus_wreq_addr,
      bus_wreq_len                             => s_Str_bus_wreq_len,
      bus_wdat_valid                           => s_Str_bus_wdat_valid,
      bus_wdat_ready                           => s_Str_bus_wdat_ready,
      bus_wdat_data                            => s_Str_bus_wdat_data,
      bus_wdat_strobe                          => s_Str_bus_wdat_strobe,
      bus_wdat_last                            => s_Str_bus_wdat_last,
      unlock_valid                             => s_Str_unl_valid,
      unlock_ready                             => s_Str_unl_ready,
      unlock_tag                               => s_Str_unl_tag
    );

  -- Controller instance.
  UserCoreController_inst: UserCoreController
    generic map (
      REG_WIDTH                                => REG_WIDTH
    )
    port map (
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      status                                   => regs_out(2*REG_WIDTH-1 downto REG_WIDTH),
      control                                  => regs_in(REG_WIDTH-1 downto 0),
      start                                    => uctrl_start,
      stop                                     => uctrl_stop,
      reset                                    => uctrl_reset,
      idle                                     => uctrl_idle,
      busy                                     => uctrl_busy,
      done                                     => uctrl_done
    );

  -- Hardware Accelerated Function instance.
  stringwrite_usercore_inst: stringwrite_usercore
    generic map (
      NUM_USER_REGS                            => NUM_USER_REGS,
      TAG_WIDTH                                => TAG_WIDTH,
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      INDEX_WIDTH                              => INDEX_WIDTH,
      REG_WIDTH                                => REG_WIDTH
    )
    port map (
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      ctrl_start                               => uctrl_start,
      ctrl_stop                                => uctrl_stop,
      ctrl_reset                               => uctrl_reset,
      ctrl_idle                                => uctrl_idle,
      ctrl_busy                                => uctrl_busy,
      ctrl_done                                => uctrl_done,
      Str_in_valid                             => s_Str_in_valid(0),
      Str_in_ready                             => s_Str_in_ready(0),
      Str_in_last                              => s_Str_in_last(0),
      Str_in_length                            => s_Str_in_data(INDEX_WIDTH-1 downto 0),
      Str_in_dvalid                            => s_Str_in_dvalid(0),
      Str_in_values_in_valid                   => s_Str_in_valid(1),
      Str_in_values_in_ready                   => s_Str_in_ready(1),
      Str_in_values_in_last                    => s_Str_in_last(1),
      Str_in_values_in_dvalid                  => s_Str_in_dvalid(1),
      Str_in_values_in_data                    => s_Str_in_data(INDEX_WIDTH+511 downto INDEX_WIDTH),
      Str_in_values_in_count                   => s_Str_in_data(INDEX_WIDTH+518 downto INDEX_WIDTH+512),
      Str_cmd_valid                            => s_Str_cmd_valid,
      Str_cmd_ready                            => s_Str_cmd_ready,
      Str_cmd_firstIdx                         => s_Str_cmd_firstIdx(INDEX_WIDTH-1 downto 0),
      Str_cmd_lastIdx                          => s_Str_cmd_lastIdx(INDEX_WIDTH-1 downto 0),
      Str_cmd_tag                              => s_Str_cmd_tag(TAG_WIDTH-1 downto 0),
      Str_cmd_Str_offsets_addr                 => s_Str_cmd_ctrl(BUS_ADDR_WIDTH-1 downto 0),
      Str_cmd_Str_values_addr                  => s_Str_cmd_ctrl(BUS_ADDR_WIDTH+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH),
      Str_unl_ready                            => s_Str_unl_ready,
      Str_unl_valid                            => s_Str_unl_valid,
      Str_unl_tag                              => s_Str_unl_tag,
      idx_first                                => regs_in(5*REG_WIDTH-1 downto 4*REG_WIDTH),
      idx_last                                 => regs_in(6*REG_WIDTH-1 downto 5*REG_WIDTH),
      reg_return0                              => regs_out(3*REG_WIDTH-1 downto 2*REG_WIDTH),
      reg_return1                              => regs_out(4*REG_WIDTH-1 downto 3*REG_WIDTH),
      reg_Str_offsets_addr                     => regs_in(8*REG_WIDTH-1 downto 6*REG_WIDTH),
      reg_Str_values_addr                      => regs_in(10*REG_WIDTH-1 downto 8*REG_WIDTH),
      regs_in                                  => s_regs_in,
      regs_out                                 => s_regs_out,
      regs_out_en                              => s_regs_out_en
    );

  -- Arbiter instance generated to serve 1 column writers.
  BusWriteArbiterVec_inst: BusWriteArbiterVec
    generic map (
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH                            => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH                           => BUS_DATA_WIDTH,
      BUS_STROBE_WIDTH                         => BUS_STROBE_WIDTH,
      NUM_SLAVE_PORTS                          => 1
    )
    port map (
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      bsv_wdat_valid                           => s_bsv_wdat_valid,
      bsv_wdat_ready                           => s_bsv_wdat_ready,
      bsv_wdat_data                            => s_bsv_wdat_data,
      bsv_wdat_strobe                          => s_bsv_wdat_strobe,
      bsv_wdat_last                            => s_bsv_wdat_last,
      bsv_wreq_valid                           => s_bsv_wreq_valid,
      bsv_wreq_ready                           => s_bsv_wreq_ready,
      bsv_wreq_addr                            => s_bsv_wreq_addr,
      bsv_wreq_len                             => s_bsv_wreq_len,
      mst_wreq_valid                           => mst_wreq_valid,
      mst_wreq_ready                           => mst_wreq_ready,
      mst_wreq_addr                            => mst_wreq_addr,
      mst_wreq_len                             => mst_wreq_len,
      mst_wdat_valid                           => mst_wdat_valid,
      mst_wdat_ready                           => mst_wdat_ready,
      mst_wdat_data                            => mst_wdat_data,
      mst_wdat_strobe                          => mst_wdat_strobe,
      mst_wdat_last                            => mst_wdat_last
    );


  regs_out(NUM_REGS*REG_WIDTH-1 downto (NUM_REGS-NUM_USER_REGS)*REG_WIDTH)<= s_regs_out;
  regs_out_en(NUM_REGS-1 downto NUM_REGS-NUM_USER_REGS)<= s_regs_out_en;
  s_regs_in                                    <= regs_in(NUM_REGS*REG_WIDTH-1 downto (NUM_REGS-NUM_USER_REGS)*REG_WIDTH);
  -----------------------------------------------------------------------------
  s_bsv_wreq_addr(BUS_ADDR_WIDTH-1 downto 0)   <= s_Str_bus_wreq_addr;
  s_bsv_wreq_len(BUS_LEN_WIDTH-1 downto 0)     <= s_Str_bus_wreq_len;
  s_Str_bus_wreq_ready                         <= s_bsv_wreq_ready(0);
  s_bsv_wreq_valid(0)                          <= s_Str_bus_wreq_valid;
  -----------------------------------------------------------------------------
  s_bsv_wdat_data(BUS_DATA_WIDTH-1 downto 0)   <= s_Str_bus_wdat_data;
  s_bsv_wdat_last(0)                           <= s_Str_bus_wdat_last;
  s_Str_bus_wdat_ready                         <= s_bsv_wdat_ready(0);
  s_bsv_wdat_strobe(BUS_STROBE_WIDTH-1 downto 0)<= s_Str_bus_wdat_strobe;
  s_bsv_wdat_valid(0)                          <= s_Str_bus_wdat_valid;
  -----------------------------------------------------------------------------
  mst_rreq_valid                               <='0';
  mst_rdat_ready                               <='0';
  regs_out_en(0)                               <='0';
  regs_out_en(1)                               <='1';
  regs_out_en(2)                               <='1';
  regs_out_en(3)                               <='1';

end architecture;

