-- Copyright 2018 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.

-- This file was automatically generated by FletchGen. Modify this file
-- at your own risk.

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

library work;
  use work.Streams.all;

entity filter_usercore is
  generic(
    TAG_WIDTH                                  : natural;
    BUS_ADDR_WIDTH                             : natural;
    INDEX_WIDTH                                : natural;
    REG_WIDTH                                  : natural
  );
  port(
    write_first_name_unlock_valid              : in std_logic;
    write_first_name_unlock_tag                : in std_logic_vector(TAG_WIDTH-1 downto 0) := (others => '0');
    write_first_name_unlock_ready              : out std_logic;
    write_first_name_in_values_in_valid        : out std_logic;
    write_first_name_in_values_in_ready        : in std_logic;
    write_first_name_in_values_in_last         : out std_logic;
    write_first_name_in_values_in_dvalid       : out std_logic;
    write_first_name_in_values_in_data         : out std_logic_vector(7 downto 0);
    write_first_name_in_values_in_count        : out std_logic_vector(0 downto 0);
    write_first_name_in_valid                  : out std_logic;
    write_first_name_in_ready                  : in std_logic;
    write_first_name_in_length                 : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    write_first_name_in_last                   : out std_logic;
    write_first_name_cmd_write_first_name_values_addr: out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    write_first_name_cmd_write_first_name_offsets_addr: out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    write_first_name_cmd_valid                 : out std_logic;
    write_first_name_cmd_tag                   : out std_logic_vector(TAG_WIDTH-1 downto 0);
    write_first_name_cmd_ready                 : in std_logic;
    write_first_name_cmd_lastIdx               : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    write_first_name_cmd_firstIdx              : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    -------------------------------------------------------------------------
    reg_write_first_name_values_addr           : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    reg_write_first_name_offsets_addr          : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    -------------------------------------------------------------------------
    reg_return1                                : out std_logic_vector(REG_WIDTH-1 downto 0);
    reg_return0                                : out std_logic_vector(REG_WIDTH-1 downto 0);
    -------------------------------------------------------------------------
    reg_read_zipcode_values_addr               : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    reg_read_last_name_values_addr             : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    reg_read_last_name_offsets_addr            : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    reg_read_first_name_values_addr            : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    reg_read_first_name_offsets_addr           : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    -------------------------------------------------------------------------
    read_zipcode_unlock_valid                  : in std_logic;
    read_zipcode_unlock_tag                    : in std_logic_vector(TAG_WIDTH-1 downto 0);
    read_zipcode_unlock_ready                  : out std_logic;
    read_zipcode_out_valid                     : in std_logic;
    read_zipcode_out_ready                     : out std_logic;
    read_zipcode_out_last                      : in std_logic;
    read_zipcode_out_data                      : in std_logic_vector(31 downto 0);
    read_zipcode_cmd_valid                     : out std_logic;
    read_zipcode_cmd_tag                       : out std_logic_vector(TAG_WIDTH-1 downto 0);
    read_zipcode_cmd_ready                     : in std_logic;
    read_zipcode_cmd_read_zipcode_values_addr  : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    read_zipcode_cmd_lastIdx                   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    read_zipcode_cmd_firstIdx                  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    read_last_name_unlock_valid                : in std_logic;
    read_last_name_unlock_tag                  : in std_logic_vector(TAG_WIDTH-1 downto 0);
    read_last_name_unlock_ready                : out std_logic;
    read_last_name_out_values_out_valid        : in std_logic;
    read_last_name_out_values_out_ready        : out std_logic;
    read_last_name_out_values_out_last         : in std_logic;
    read_last_name_out_values_out_dvalid       : in std_logic;
    read_last_name_out_values_out_data         : in std_logic_vector(7 downto 0);
    read_last_name_out_values_out_count        : in std_logic_vector(0 downto 0);
    read_last_name_out_valid                   : in std_logic;
    read_last_name_out_ready                   : out std_logic;
    read_last_name_out_length                  : in std_logic_vector(INDEX_WIDTH-1 downto 0);
    read_last_name_out_last                    : in std_logic;
    read_last_name_cmd_valid                   : out std_logic;
    read_last_name_cmd_tag                     : out std_logic_vector(TAG_WIDTH-1 downto 0);
    read_last_name_cmd_ready                   : in std_logic;
    read_last_name_cmd_read_last_name_values_addr: out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    read_last_name_cmd_read_last_name_offsets_addr: out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    read_last_name_cmd_lastIdx                 : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    read_last_name_cmd_firstIdx                : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    read_first_name_unlock_valid               : in std_logic;
    read_first_name_unlock_tag                 : in std_logic_vector(TAG_WIDTH-1 downto 0);
    read_first_name_unlock_ready               : out std_logic;
    read_first_name_out_values_out_valid       : in std_logic;
    read_first_name_out_values_out_ready       : out std_logic;
    read_first_name_out_values_out_last        : in std_logic;
    read_first_name_out_values_out_dvalid      : in std_logic;
    read_first_name_out_values_out_data        : in std_logic_vector(7 downto 0);
    read_first_name_out_values_out_count       : in std_logic_vector(0 downto 0);
    read_first_name_out_valid                  : in std_logic;
    read_first_name_out_ready                  : out std_logic;
    read_first_name_out_length                 : in std_logic_vector(INDEX_WIDTH-1 downto 0);
    read_first_name_out_last                   : in std_logic;
    read_first_name_cmd_valid                  : out std_logic;
    read_first_name_cmd_tag                    : out std_logic_vector(TAG_WIDTH-1 downto 0);
    read_first_name_cmd_ready                  : in std_logic;
    read_first_name_cmd_read_first_name_values_addr: out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    read_first_name_cmd_read_first_name_offsets_addr: out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    read_first_name_cmd_lastIdx                : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    read_first_name_cmd_firstIdx               : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    -------------------------------------------------------------------------
    idx_last                                   : in std_logic_vector(REG_WIDTH-1 downto 0);
    idx_first                                  : in std_logic_vector(REG_WIDTH-1 downto 0);
    -------------------------------------------------------------------------
    ctrl_stop                                  : in std_logic;
    ctrl_start                                 : in std_logic;
    ctrl_reset                                 : in std_logic;
    ctrl_idle                                  : out std_logic;
    ctrl_done                                  : out std_logic;
    ctrl_busy                                  : out std_logic;
    -------------------------------------------------------------------------
    acc_reset                                  : in std_logic;
    acc_clk                                    : in std_logic
  );
end entity;

architecture Implementation of filter_usercore is

  component filter_hls_fletcher is
  port (
      ap_clk : IN STD_LOGIC;
      ap_rst : IN STD_LOGIC;
      ap_start : IN STD_LOGIC;
      ap_done : OUT STD_LOGIC;
      ap_idle : OUT STD_LOGIC;
      ap_ready : OUT STD_LOGIC;
      num_entries : IN STD_LOGIC_VECTOR (31 downto 0);
      in_first_name_length_V_dout : IN STD_LOGIC_VECTOR (31 downto 0);
      in_first_name_length_V_empty_n : IN STD_LOGIC;
      in_first_name_length_V_read : OUT STD_LOGIC;
      in_first_name_values_V_dout : IN STD_LOGIC_VECTOR (7 downto 0);
      in_first_name_values_V_empty_n : IN STD_LOGIC;
      in_first_name_values_V_read : OUT STD_LOGIC;
      in_last_name_length_V_dout : IN STD_LOGIC_VECTOR (31 downto 0);
      in_last_name_length_V_empty_n : IN STD_LOGIC;
      in_last_name_length_V_read : OUT STD_LOGIC;
      in_last_name_values_V_dout : IN STD_LOGIC_VECTOR (7 downto 0);
      in_last_name_values_V_empty_n : IN STD_LOGIC;
      in_last_name_values_V_read : OUT STD_LOGIC;
      in_zipcode_V_dout : IN STD_LOGIC_VECTOR (31 downto 0);
      in_zipcode_V_empty_n : IN STD_LOGIC;
      in_zipcode_V_read : OUT STD_LOGIC;
      filter_name_address0 : OUT STD_LOGIC_VECTOR (5 downto 0);
      filter_name_ce0 : OUT STD_LOGIC;
      filter_name_q0 : IN STD_LOGIC_VECTOR (7 downto 0);
      filter_zipcode : IN STD_LOGIC_VECTOR (31 downto 0);
      out_first_name_length_V_din : OUT STD_LOGIC_VECTOR (31 downto 0);
      out_first_name_length_V_full_n : IN STD_LOGIC;
      out_first_name_length_V_write : OUT STD_LOGIC;
      out_first_name_values_V_din : OUT STD_LOGIC_VECTOR (7 downto 0);
      out_first_name_values_V_full_n : IN STD_LOGIC;
      out_first_name_values_V_write : OUT STD_LOGIC;
      ap_return : OUT STD_LOGIC_VECTOR (31 downto 0));
  end component;

  type read_cmd_type is record
    valid                     : std_logic;
    ready                     : std_logic;
    tag                       : std_logic_vector(TAG_WIDTH-1 downto 0);
    lastIdx                   : std_logic_vector(INDEX_WIDTH-1 downto 0);
    firstIdx                  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  end record;
  
  type write_cmd_type is record
    valid                     : std_logic;
    ready                     : std_logic;
    tag                       : std_logic_vector(TAG_WIDTH-1 downto 0);
    lastIdx                   : std_logic_vector(INDEX_WIDTH-1 downto 0);
    firstIdx                  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  end record;

  type unlock_type is record
    valid                     : std_logic;
    ready                     : std_logic;
  end record;

  type hls_cin_type is record
    start             : std_logic;
    reset             : std_logic;
  end record;

  type hls_cout_type is record
    idle              : std_logic;
    done              : std_logic;
    ready             : std_logic;
  end record;

  type hls_arg_type is record
    num_entries       : std_logic_vector (31 downto 0);
    filter_zipcode    : std_logic_vector (31 downto 0);
  end record;
  
  type hls_ret_type is record
    ret               : std_logic_vector(31 downto 0);
  end record;

  type hls_din_type is record
    fn_length_data     : STD_LOGIC_VECTOR (31 downto 0);
    fn_length_valid    : STD_LOGIC;
    fn_length_ready    : STD_LOGIC;
    fn_values_data     : STD_LOGIC_VECTOR (7 downto 0);
    fn_values_valid    : STD_LOGIC;
    fn_values_ready    : STD_LOGIC;
    ln_length_data     : STD_LOGIC_VECTOR (31 downto 0);
    ln_length_valid    : STD_LOGIC;
    ln_length_ready    : STD_LOGIC;
    ln_values_data     : STD_LOGIC_VECTOR (7 downto 0);
    ln_values_valid    : STD_LOGIC;
    ln_values_ready    : STD_LOGIC;
    zip_data           : STD_LOGIC_VECTOR (31 downto 0);
    zip_valid          : STD_LOGIC;
    zip_ready          : STD_LOGIC;
  end record;

  type hls_dout_type is record
    fn_length_data     : STD_LOGIC_VECTOR (31 downto 0);
    fn_length_valid    : STD_LOGIC;
    fn_length_ready    : STD_LOGIC;
    fn_values_data     : STD_LOGIC_VECTOR (7 downto 0);
    fn_values_valid    : STD_LOGIC;
    fn_values_ready    : STD_LOGIC;
  end record;

  type hls_name_type is record
    addr              : STD_LOGIC_VECTOR (5 downto 0);
    ce                : STD_LOGIC;
    q                 : STD_LOGIC_VECTOR (7 downto 0);
  end record;


  type state_type is (IDLE, RD_CMD, WR_CMD, BUSY, FINISH_VAL, FINISH_LEN, UNL, DONE);

  type reg_record is record
    busy                      : std_logic;
    done                      : std_logic;
    reset_start               : std_logic;
    state                     : state_type;
  end record;

  signal r : reg_record;
  signal d : reg_record;
  
  signal read_cmd               : read_cmd_type;
  signal write_cmd              : write_cmd_type;
  signal unlock                 : unlock_type;

  signal hls_cin                : hls_cin_type;
  signal hls_args               : hls_arg_type;
  signal hls_name               : hls_name_type;
  signal hls_din                : hls_din_type;
  signal hls_cout               : hls_cout_type;
  signal hls_ret                : hls_ret_type;
  signal hls_dout               : hls_dout_type;
  
  type name_ram_type is array (63 downto 0) of Character;
  
  signal name_ram : name_ram_type := (
    0 => 'S',
    1 => 'm',
    2 => 'i',
    3 => 't',
    4 => 'h',
    others => nul
  );

begin
  -- Connect all addresses
  read_zipcode_cmd_read_zipcode_values_addr          <= reg_read_zipcode_values_addr;
  read_last_name_cmd_read_last_name_values_addr      <= reg_read_last_name_values_addr;
  read_last_name_cmd_read_last_name_offsets_addr     <= reg_read_last_name_offsets_addr;
  read_first_name_cmd_read_first_name_values_addr    <= reg_read_first_name_values_addr;
  read_first_name_cmd_read_first_name_offsets_addr   <= reg_read_first_name_offsets_addr;
  write_first_name_cmd_write_first_name_values_addr  <= reg_write_first_name_values_addr;
  write_first_name_cmd_write_first_name_offsets_addr <= reg_write_first_name_offsets_addr;

  -- Get first and last idx from registers
  read_cmd.firstIdx  <= idx_first;
  read_cmd.lastIdx   <= idx_last;
  
  -- We don't know howmany entries will match the filter so 
  -- set both first and last index to 0.
  write_cmd.firstIdx <= (others => '0');
  write_cmd.lastIdx  <= (others => '0');

  read_cmd.tag                  <= (others => '0');
  write_cmd.tag                 <= (others => '0');

  -- Connect all command streams, combine read commands
  read_first_name_cmd_tag       <= read_cmd.tag;
  read_last_name_cmd_tag        <= read_cmd.tag;
  read_zipcode_cmd_tag          <= read_cmd.tag;
  write_first_name_cmd_tag      <= write_cmd.tag;

  read_first_name_cmd_firstIdx  <= read_cmd.firstIdx;
  read_last_name_cmd_firstIdx   <= read_cmd.firstIdx;
  read_zipcode_cmd_firstIdx     <= read_cmd.firstIdx;
  write_first_name_cmd_firstIdx <= write_cmd.firstIdx;

  read_first_name_cmd_lastIdx   <= read_cmd.lastIdx;
  read_last_name_cmd_lastIdx    <= read_cmd.lastIdx;
  read_zipcode_cmd_lastIdx      <= read_cmd.lastIdx;
  write_first_name_cmd_lastIdx  <= write_cmd.lastIdx;

  -- Synchronize the three command streams from the input columns
  read_cmd_sync : StreamSync
    generic map (
      NUM_INPUTS => 1,
      NUM_OUTPUTS => 3
    )
    port map (
      clk   => acc_clk,
      reset => acc_reset,
      in_valid(0) => read_cmd.valid,
      in_ready(0) => read_cmd.ready,
      out_valid(0) => read_first_name_cmd_valid,
      out_valid(1) => read_last_name_cmd_valid,
      out_valid(2) => read_zipcode_cmd_valid,
      out_ready(0) => read_first_name_cmd_ready,
      out_ready(1) => read_last_name_cmd_ready,
      out_ready(2) => read_zipcode_cmd_ready
    );
    
  write_first_name_cmd_valid <= write_cmd.valid;
  write_cmd.ready <= write_first_name_cmd_ready;

  -- Synchronize the four unlock streams
  read_unlock_sync : StreamSync
    generic map (
      NUM_INPUTS => 3,
      NUM_OUTPUTS => 1
    )
    port map (
      clk   => acc_clk,
      reset => acc_reset,
      in_valid(0) => read_first_name_unlock_valid,
      in_valid(1) => read_last_name_unlock_valid,
      in_valid(2) => read_zipcode_unlock_valid,
      in_ready(0) => read_first_name_unlock_ready,
      in_ready(1) => read_last_name_unlock_ready,
      in_ready(2) => read_zipcode_unlock_ready,
      
      out_valid(0) => unlock.valid,
      out_ready(0) => unlock.ready
    );
      
  read_first_name_unlock_ready  <= unlock.ready;
  read_last_name_unlock_ready   <= unlock.ready;
  read_zipcode_unlock_ready     <= unlock.ready;


  seq_proc: process(acc_clk) is
  begin
    if rising_edge(acc_clk) then
      r <= d;

      -- Reset
      if acc_reset = '1' then
        r.state         <= IDLE;
        r.reset_start   <= '0';
        r.busy          <= '0';
        r.done          <= '0';
      end if;
    end if;
  end process;

  comb_proc: process(all) is
    variable v : reg_record;
  begin
    -- Default registered outputs:
    v := r;

    -- Default combinatorial outputs:
    read_cmd.valid  <= '0';
    write_cmd.valid <= '0';
    unlock.ready    <= '0';
    
    write_first_name_unlock_ready        <= '0';
    
    write_first_name_in_values_in_data   <= (others => '1');
    write_first_name_in_values_in_last   <= '0';
    write_first_name_in_values_in_dvalid <= '0';
    write_first_name_in_values_in_valid  <= '0';
    
    write_first_name_in_length           <= (others => '0'); 
    write_first_name_in_last             <= '0';
    write_first_name_in_valid            <= '0';
    
    hls_args.num_entries <= idx_last;
    hls_args.filter_zipcode <= X"00000539"; -- 1337

    case r.state is
      when IDLE =>
        ctrl_idle      <= '1';
        ctrl_busy      <= '0';
        ctrl_done      <= '0';
        hls_cin.reset  <= '1';
        hls_cin.start  <= '0';

        if ctrl_start = '1' then
          v.reset_start := '1';
          v.state := RD_CMD;
          v.busy := '1';
          v.done := '0';
        end if;
        
      when RD_CMD =>
        ctrl_idle      <= '0';
        ctrl_busy      <= '1';
        ctrl_done      <= '0';
        hls_cin.reset  <= '0';
        hls_cin.start  <= '1';

        read_cmd.valid <= '1';
        if read_cmd.ready = '1' then
          v.state := WR_CMD;
        end if;
        
      when WR_CMD =>
        ctrl_idle      <= '0';
        ctrl_busy      <= '1';
        ctrl_done      <= '0';
        hls_cin.reset  <= '0';
        hls_cin.start  <= '0';       
        
        write_cmd.valid <= '1';
        if (write_cmd.ready = '1') then
          v.state := BUSY;
        end if;        
        
      when BUSY =>
        ctrl_idle      <= '0';
        ctrl_busy      <= '1';
        ctrl_done      <= '0';
        hls_cin.reset  <= '0';
        hls_cin.start  <= '0';
       
       -- Pass-through the data
        write_first_name_in_values_in_last   <= '0';
        write_first_name_in_values_in_dvalid <= '1';
        write_first_name_in_values_in_valid  <= hls_dout.fn_values_valid;
        write_first_name_in_values_in_data   <= hls_dout.fn_values_data;
        write_first_name_in_valid            <= hls_dout.fn_length_valid;
        write_first_name_in_length           <= hls_dout.fn_length_data; 
        write_first_name_in_last             <= '0';       
        
        if unlock.valid = '1' and
           hls_cout.done = '1' and
           hls_cout.ready = '1'
        then
          unlock.ready <= '1';
          v.state := FINISH_VAL;
        end if;
        
      when FINISH_VAL =>
        ctrl_idle      <= '0';
        ctrl_busy      <= '1';
        ctrl_done      <= '0';
        hls_cin.reset  <= '0';
        hls_cin.start  <= '0';
       
        -- Create a handshake 
        write_first_name_in_values_in_last   <= '1';
        write_first_name_in_values_in_valid  <= '1';
        
        if write_first_name_in_values_in_ready <= '1' then
           v.state := FINISH_LEN;
        end if;

      when FINISH_LEN =>
        ctrl_idle      <= '0';
        ctrl_busy      <= '1';
        ctrl_done      <= '0';
        hls_cin.reset  <= '0';
        hls_cin.start  <= '0';
        
        write_first_name_in_valid            <= '1';
        write_first_name_in_last             <= '1';
        
        if write_first_name_in_ready = '1' then
           v.state := UNL;
        end if;
        
      when UNL =>
        ctrl_idle      <= '0';
        ctrl_busy      <= '1';
        ctrl_done      <= '0';
        hls_cin.reset  <= '0';
        hls_cin.start  <= '0';
        
        if write_first_name_unlock_valid = '1' then
          write_first_name_unlock_ready <= '1';
          v.state := DONE;
        end if;
        
      when DONE =>
        ctrl_idle      <= '0';
        ctrl_busy      <= '0';
        ctrl_done      <= '1';
        hls_cin.reset  <= '0';
        hls_cin.start  <= '0';

    end case;

    d <= v;

  end process;

  hls_core: filter_hls_fletcher
    port map (
        ap_clk                            => acc_clk,
        ap_rst                            => hls_cin.reset,
        ap_start                          => hls_cin.start,
        ap_done                           => hls_cout.done,
        ap_idle                           => hls_cout.idle,
        ap_ready                          => hls_cout.ready,
        num_entries                       => hls_args.num_entries,
        in_first_name_length_V_dout       => hls_din.fn_length_data,
        in_first_name_length_V_empty_n    => hls_din.fn_length_valid,
        in_first_name_length_V_read       => hls_din.fn_length_ready,
        in_first_name_values_V_dout       => hls_din.fn_values_data,
        in_first_name_values_V_empty_n    => hls_din.fn_values_valid,
        in_first_name_values_V_read       => hls_din.fn_values_ready,
        in_last_name_length_V_dout        => hls_din.ln_length_data,
        in_last_name_length_V_empty_n     => hls_din.ln_length_valid,
        in_last_name_length_V_read        => hls_din.ln_length_ready,
        in_last_name_values_V_dout        => hls_din.ln_values_data,
        in_last_name_values_V_empty_n     => hls_din.ln_values_valid,
        in_last_name_values_V_read        => hls_din.ln_values_ready,
        in_zipcode_V_dout                 => hls_din.zip_data,
        in_zipcode_V_empty_n              => hls_din.zip_valid,
        in_zipcode_V_read                 => hls_din.zip_ready,
        filter_name_address0              => hls_name.addr,
        filter_name_ce0                   => hls_name.ce,
        filter_name_q0                    => hls_name.q,
        filter_zipcode                    => hls_args.filter_zipcode,
        out_first_name_length_V_din       => hls_dout.fn_length_data,
        out_first_name_length_V_full_n    => hls_dout.fn_length_ready,
        out_first_name_length_V_write     => hls_dout.fn_length_valid,
        out_first_name_values_V_din       => hls_dout.fn_values_data,
        out_first_name_values_V_full_n    => hls_dout.fn_values_ready,
        out_first_name_values_V_write     => hls_dout.fn_values_valid,
        ap_return                         => hls_ret.ret
    );

    -- HLS core input streams
    hls_din.fn_length_data                <= read_first_name_out_length;
    hls_din.fn_length_valid               <= read_first_name_out_valid;
    read_last_name_out_ready              <= hls_din.fn_length_ready;
    hls_din.fn_values_data                <= read_first_name_out_values_out_data;
    hls_din.fn_values_valid               <= read_first_name_out_values_out_valid;
    read_first_name_out_values_out_ready  <= hls_din.fn_values_ready;
    hls_din.ln_length_data                <= read_last_name_out_length;
    hls_din.ln_length_valid               <= read_last_name_out_valid;
    read_first_name_out_ready             <= hls_din.ln_length_ready;
    hls_din.ln_values_data                <= read_last_name_out_values_out_data;
    hls_din.ln_values_valid               <= read_last_name_out_values_out_valid;
    read_last_name_out_values_out_ready   <= hls_din.ln_values_ready;
    hls_din.zip_data                      <= read_zipcode_out_data;
    hls_din.zip_valid                     <= read_zipcode_out_valid;
    read_zipcode_out_ready                <= hls_din.zip_ready;
    
    -- HLS core output streams
    hls_dout.fn_length_ready              <= write_first_name_in_ready;
    hls_dout.fn_values_ready              <= write_first_name_in_values_in_ready;

    -- filter name parameter RAM
    name_ram_proc: process(acc_clk) is
    begin
      if rising_edge(acc_clk) then
        if hls_name.ce = '1' then
          hls_name.q <= std_logic_vector(to_unsigned(character'pos(name_ram(to_integer(unsigned(hls_name.addr)))),8));
        end if;
      end if;
    end process;
    

end architecture;
