-- Copyright 2018 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.

-- This file was automatically generated by FletchGen. Modify this file
-- at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;

library work;
use work.Arrow.all;
use work.Arrays.all;
use work.Interconnect.all;
use work.Wrapper.all;

entity filter_wrapper is
  generic(
    BUS_ADDR_WIDTH                             : natural;
    BUS_DATA_WIDTH                             : natural;
    BUS_STROBE_WIDTH                           : natural;
    BUS_LEN_WIDTH                              : natural;
    BUS_BURST_STEP_LEN                         : natural;
    BUS_BURST_MAX_LEN                          : natural;
    ---------------------------------------------------------------------------
    INDEX_WIDTH                                : natural;
    ---------------------------------------------------------------------------
    NUM_ARROW_BUFFERS                          : natural;
    NUM_REGS                                   : natural;
    NUM_USER_REGS                              : natural;
    REG_WIDTH                                  : natural;
    ---------------------------------------------------------------------------
    TAG_WIDTH                                  : natural
  );
  port(
    acc_reset                                  : in std_logic;
    bus_clk                                    : in std_logic;
    bus_reset                                  : in std_logic;
    acc_clk                                    : in std_logic;
    ---------------------------------------------------------------------------
    mst_rreq_valid                             : out std_logic;
    mst_rreq_ready                             : in std_logic;
    mst_rreq_addr                              : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    mst_rreq_len                               : out std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
    ---------------------------------------------------------------------------
    mst_rdat_valid                             : in std_logic;
    mst_rdat_ready                             : out std_logic;
    mst_rdat_data                              : in std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
    mst_rdat_last                              : in std_logic;
    ---------------------------------------------------------------------------
    mst_wreq_valid                             : out std_logic;
    mst_wreq_len                               : out std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
    mst_wreq_addr                              : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    mst_wreq_ready                             : in std_logic;
    ---------------------------------------------------------------------------
    mst_wdat_valid                             : out std_logic;
    mst_wdat_ready                             : in std_logic;
    mst_wdat_data                              : out std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
    mst_wdat_strobe                            : out std_logic_vector(BUS_STROBE_WIDTH-1 downto 0);
    mst_wdat_last                              : out std_logic;
    ---------------------------------------------------------------------------
    regs_in                                    : in std_logic_vector(NUM_REGS*REG_WIDTH-1 downto 0);
    regs_out                                   : out std_logic_vector(NUM_REGS*REG_WIDTH-1 downto 0);
    regs_out_en                                : out std_logic_vector(NUM_REGS-1 downto 0)
  );
end filter_wrapper;

architecture Implementation of filter_wrapper is

  -----------------------------------------------------------------------------
  -- Hardware Accelerated Function component.
  -- This component should be implemented by the user.
  component filter_usercore is
    generic(
      TAG_WIDTH                                  : natural;
      BUS_ADDR_WIDTH                             : natural;
      INDEX_WIDTH                                : natural;
      REG_WIDTH                                  : natural
    );
    port(
      write_first_name_unlock_valid              : in std_logic;
      write_first_name_unlock_tag                : in std_logic_vector(TAG_WIDTH-1 downto 0);
      write_first_name_unlock_ready              : out std_logic;
      write_first_name_in_values_in_valid        : out std_logic;
      write_first_name_in_values_in_ready        : in std_logic;
      write_first_name_in_values_in_last         : out std_logic;
      write_first_name_in_values_in_dvalid       : out std_logic;
      write_first_name_in_values_in_data         : out std_logic_vector(7 downto 0);
      write_first_name_in_values_in_count        : out std_logic_vector(0 downto 0);
      write_first_name_in_valid                  : out std_logic;
      write_first_name_in_ready                  : in std_logic;
      write_first_name_in_length                 : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      write_first_name_in_last                   : out std_logic;
      write_first_name_cmd_write_first_name_values_addr: out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      write_first_name_cmd_write_first_name_offsets_addr: out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      write_first_name_cmd_valid                 : out std_logic;
      write_first_name_cmd_tag                   : out std_logic_vector(TAG_WIDTH-1 downto 0);
      write_first_name_cmd_ready                 : in std_logic;
      write_first_name_cmd_lastIdx               : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      write_first_name_cmd_firstIdx              : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      -------------------------------------------------------------------------
      reg_write_first_name_values_addr           : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      reg_write_first_name_offsets_addr          : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      -------------------------------------------------------------------------
      reg_return1                                : out std_logic_vector(REG_WIDTH-1 downto 0);
      reg_return0                                : out std_logic_vector(REG_WIDTH-1 downto 0);
      -------------------------------------------------------------------------
      reg_read_zipcode_values_addr               : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      reg_read_last_name_values_addr             : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      reg_read_last_name_offsets_addr            : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      reg_read_first_name_values_addr            : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      reg_read_first_name_offsets_addr           : in std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      -------------------------------------------------------------------------
      read_zipcode_unlock_valid                  : in std_logic;
      read_zipcode_unlock_tag                    : in std_logic_vector(TAG_WIDTH-1 downto 0);
      read_zipcode_unlock_ready                  : out std_logic;
      read_zipcode_out_valid                     : in std_logic;
      read_zipcode_out_ready                     : out std_logic;
      read_zipcode_out_last                      : in std_logic;
      read_zipcode_out_data                      : in std_logic_vector(31 downto 0);
      read_zipcode_cmd_valid                     : out std_logic;
      read_zipcode_cmd_tag                       : out std_logic_vector(TAG_WIDTH-1 downto 0);
      read_zipcode_cmd_ready                     : in std_logic;
      read_zipcode_cmd_read_zipcode_values_addr  : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      read_zipcode_cmd_lastIdx                   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      read_zipcode_cmd_firstIdx                  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      read_last_name_unlock_valid                : in std_logic;
      read_last_name_unlock_tag                  : in std_logic_vector(TAG_WIDTH-1 downto 0);
      read_last_name_unlock_ready                : out std_logic;
      read_last_name_out_values_out_valid        : in std_logic;
      read_last_name_out_values_out_ready        : out std_logic;
      read_last_name_out_values_out_last         : in std_logic;
      read_last_name_out_values_out_dvalid       : in std_logic;
      read_last_name_out_values_out_data         : in std_logic_vector(7 downto 0);
      read_last_name_out_values_out_count        : in std_logic_vector(0 downto 0);
      read_last_name_out_valid                   : in std_logic;
      read_last_name_out_ready                   : out std_logic;
      read_last_name_out_length                  : in std_logic_vector(INDEX_WIDTH-1 downto 0);
      read_last_name_out_last                    : in std_logic;
      read_last_name_cmd_valid                   : out std_logic;
      read_last_name_cmd_tag                     : out std_logic_vector(TAG_WIDTH-1 downto 0);
      read_last_name_cmd_ready                   : in std_logic;
      read_last_name_cmd_read_last_name_values_addr: out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      read_last_name_cmd_read_last_name_offsets_addr: out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      read_last_name_cmd_lastIdx                 : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      read_last_name_cmd_firstIdx                : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      read_first_name_unlock_valid               : in std_logic;
      read_first_name_unlock_tag                 : in std_logic_vector(TAG_WIDTH-1 downto 0);
      read_first_name_unlock_ready               : out std_logic;
      read_first_name_out_values_out_valid       : in std_logic;
      read_first_name_out_values_out_ready       : out std_logic;
      read_first_name_out_values_out_last        : in std_logic;
      read_first_name_out_values_out_dvalid      : in std_logic;
      read_first_name_out_values_out_data        : in std_logic_vector(7 downto 0);
      read_first_name_out_values_out_count       : in std_logic_vector(0 downto 0);
      read_first_name_out_valid                  : in std_logic;
      read_first_name_out_ready                  : out std_logic;
      read_first_name_out_length                 : in std_logic_vector(INDEX_WIDTH-1 downto 0);
      read_first_name_out_last                   : in std_logic;
      read_first_name_cmd_valid                  : out std_logic;
      read_first_name_cmd_tag                    : out std_logic_vector(TAG_WIDTH-1 downto 0);
      read_first_name_cmd_ready                  : in std_logic;
      read_first_name_cmd_read_first_name_values_addr: out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      read_first_name_cmd_read_first_name_offsets_addr: out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
      read_first_name_cmd_lastIdx                : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      read_first_name_cmd_firstIdx               : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      -------------------------------------------------------------------------
      idx_last                                   : in std_logic_vector(REG_WIDTH-1 downto 0);
      idx_first                                  : in std_logic_vector(REG_WIDTH-1 downto 0);
      -------------------------------------------------------------------------
      ctrl_stop                                  : in std_logic;
      ctrl_start                                 : in std_logic;
      ctrl_reset                                 : in std_logic;
      ctrl_idle                                  : out std_logic;
      ctrl_done                                  : out std_logic;
      ctrl_busy                                  : out std_logic;
      -------------------------------------------------------------------------
      acc_reset                                  : in std_logic;
      acc_clk                                    : in std_logic
    );
  end component;
  -----------------------------------------------------------------------------

  signal s_read_first_name_cmd_ready           : std_logic;
  signal uctrl_done                            : std_logic;
  signal uctrl_busy                            : std_logic;
  signal uctrl_idle                            : std_logic;
  signal uctrl_reset                           : std_logic;
  signal uctrl_stop                            : std_logic;
  signal uctrl_start                           : std_logic;
  signal uctrl_control                         : std_logic_vector(REG_WIDTH-1 downto 0);
  signal uctrl_status                          : std_logic_vector(REG_WIDTH-1 downto 0);
  signal s_read_first_name_bus_rdat_last       : std_logic;
  signal s_read_first_name_bus_rdat_data       : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal s_read_first_name_bus_rdat_ready      : std_logic;
  signal s_read_first_name_bus_rdat_valid      : std_logic;
  signal s_read_first_name_bus_rreq_len        : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal s_read_first_name_bus_rreq_addr       : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_read_first_name_bus_rreq_valid      : std_logic;
  signal s_read_first_name_cmd_valid           : std_logic;
  signal s_read_first_name_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_read_first_name_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_read_first_name_cmd_ctrl            : std_logic_vector(2*BUS_ADDR_WIDTH-1 downto 0);
  signal s_read_first_name_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);
  signal s_read_first_name_unlock_valid        : std_logic;
  signal s_read_first_name_unlock_ready        : std_logic;
  signal s_read_first_name_unlock_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);
  signal s_read_first_name_bus_rreq_ready      : std_logic;
  signal s_read_first_name_out_dvalid          : std_logic_vector(1 downto 0);
  signal s_read_first_name_out_data            : std_logic_vector(INDEX_WIDTH+8 downto 0);
  signal s_read_first_name_out_last            : std_logic_vector(1 downto 0);
  signal s_read_first_name_out_ready           : std_logic_vector(1 downto 0);
  signal s_read_first_name_out_valid           : std_logic_vector(1 downto 0);
  -----------------------------------------------------------------------------
  signal s_read_last_name_cmd_lastIdx          : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_read_last_name_cmd_valid            : std_logic;
  signal s_read_last_name_cmd_ready            : std_logic;
  signal s_read_last_name_bus_rdat_last        : std_logic;
  signal s_read_last_name_bus_rdat_data        : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal s_read_last_name_bus_rdat_ready       : std_logic;
  signal s_read_last_name_bus_rdat_valid       : std_logic;
  signal s_read_last_name_bus_rreq_len         : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal s_read_last_name_bus_rreq_ready       : std_logic;
  signal s_read_last_name_cmd_firstIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_read_last_name_cmd_ctrl             : std_logic_vector(2*BUS_ADDR_WIDTH-1 downto 0);
  signal s_read_last_name_cmd_tag              : std_logic_vector(TAG_WIDTH-1 downto 0);
  signal s_read_last_name_unlock_valid         : std_logic;
  signal s_read_last_name_unlock_ready         : std_logic;
  signal s_read_last_name_unlock_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);
  signal s_read_last_name_out_valid            : std_logic_vector(1 downto 0);
  signal s_read_last_name_out_ready            : std_logic_vector(1 downto 0);
  signal s_read_last_name_bus_rreq_addr        : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_read_last_name_bus_rreq_valid       : std_logic;
  signal s_read_last_name_out_dvalid           : std_logic_vector(1 downto 0);
  signal s_read_last_name_out_data             : std_logic_vector(INDEX_WIDTH+8 downto 0);
  signal s_read_last_name_out_last             : std_logic_vector(1 downto 0);
  -----------------------------------------------------------------------------
  signal s_read_zipcode_cmd_ctrl               : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_read_zipcode_cmd_valid              : std_logic;
  signal s_read_zipcode_cmd_ready              : std_logic;
  signal s_read_zipcode_cmd_firstIdx           : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_read_zipcode_bus_rdat_last          : std_logic;
  signal s_read_zipcode_bus_rdat_data          : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal s_read_zipcode_bus_rdat_ready         : std_logic;
  signal s_read_zipcode_bus_rdat_valid         : std_logic;
  signal s_read_zipcode_bus_rreq_len           : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal s_read_zipcode_bus_rreq_ready         : std_logic;
  signal s_read_zipcode_cmd_lastIdx            : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_read_zipcode_cmd_tag                : std_logic_vector(TAG_WIDTH-1 downto 0);
  signal s_read_zipcode_unlock_valid           : std_logic;
  signal s_read_zipcode_unlock_ready           : std_logic;
  signal s_read_zipcode_unlock_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);
  signal s_read_zipcode_out_valid              : std_logic_vector(0 downto 0);
  signal s_read_zipcode_out_ready              : std_logic_vector(0 downto 0);
  signal s_read_zipcode_out_last               : std_logic_vector(0 downto 0);
  signal s_read_zipcode_bus_rreq_addr          : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_read_zipcode_bus_rreq_valid         : std_logic;
  signal s_read_zipcode_out_dvalid             : std_logic_vector(0 downto 0);
  signal s_read_zipcode_out_data               : std_logic_vector(31 downto 0);
  -----------------------------------------------------------------------------
  signal s_write_first_name_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);
  signal s_write_first_name_cmd_valid          : std_logic;
  signal s_write_first_name_cmd_ready          : std_logic;
  signal s_write_first_name_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_write_first_name_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal s_write_first_name_bus_wdat_last      : std_logic;
  signal s_write_first_name_bus_wdat_strobe    : std_logic_vector(BUS_STROBE_WIDTH-1 downto 0);
  signal s_write_first_name_bus_wdat_data      : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal s_write_first_name_bus_wdat_ready     : std_logic;
  signal s_write_first_name_bus_wdat_valid     : std_logic;
  signal s_write_first_name_bus_wreq_addr      : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_write_first_name_cmd_ctrl           : std_logic_vector(2*BUS_ADDR_WIDTH-1 downto 0);
  signal s_write_first_name_unlock_valid       : std_logic;
  signal s_write_first_name_unlock_ready       : std_logic;
  signal s_write_first_name_unlock_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);
  signal s_write_first_name_in_valid           : std_logic_vector(1 downto 0);
  signal s_write_first_name_in_ready           : std_logic_vector(1 downto 0);
  signal s_write_first_name_in_last            : std_logic_vector(1 downto 0);
  signal s_write_first_name_in_data            : std_logic_vector(INDEX_WIDTH+8 downto 0);
  signal s_write_first_name_bus_wreq_len       : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal s_write_first_name_bus_wreq_ready     : std_logic;
  signal s_write_first_name_bus_wreq_valid     : std_logic;
  signal s_write_first_name_in_dvalid          : std_logic_vector(1 downto 0);
  -----------------------------------------------------------------------------
  signal s_bsv_rreq_valid                      : std_logic_vector(2 downto 0);
  signal s_bsv_rreq_ready                      : std_logic_vector(2 downto 0);
  signal s_bsv_rreq_addr                       : std_logic_vector(3*BUS_ADDR_WIDTH-1 downto 0);
  signal s_bsv_rreq_len                        : std_logic_vector(3*BUS_LEN_WIDTH-1 downto 0);
  -----------------------------------------------------------------------------
  signal s_bsv_rdat_ready                      : std_logic_vector(2 downto 0);
  signal s_bsv_rdat_last                       : std_logic_vector(2 downto 0);
  signal s_bsv_rdat_data                       : std_logic_vector(3*BUS_DATA_WIDTH-1 downto 0);
  signal s_bsv_rdat_valid                      : std_logic_vector(2 downto 0);
  -----------------------------------------------------------------------------
  signal s_bsv_wreq_len                        : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal s_bsv_wreq_addr                       : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal s_bsv_wreq_ready                      : std_logic_vector(0 downto 0);
  signal s_bsv_wreq_valid                      : std_logic_vector(0 downto 0);
  -----------------------------------------------------------------------------
  signal s_bsv_wdat_ready                      : std_logic_vector(0 downto 0);
  signal s_bsv_wdat_data                       : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal s_bsv_wdat_strobe                     : std_logic_vector(BUS_STROBE_WIDTH-1 downto 0);
  signal s_bsv_wdat_last                       : std_logic_vector(0 downto 0);
  signal s_bsv_wdat_valid                      : std_logic_vector(0 downto 0);
begin
  -- ArrayReader instance generated from Arrow schema field:
  -- read_first_name: string not null
  read_first_name_read_inst: ArrayReader
    generic map (
      CFG                                      => "listprim(8)",
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH                            => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH                           => BUS_DATA_WIDTH,
      BUS_BURST_STEP_LEN                       => BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN                        => BUS_BURST_MAX_LEN,
      INDEX_WIDTH                              => INDEX_WIDTH,
      CMD_TAG_ENABLE                           => true
    )
    port map (
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      cmd_valid                                => s_read_first_name_cmd_valid,
      cmd_ready                                => s_read_first_name_cmd_ready,
      cmd_firstIdx                             => s_read_first_name_cmd_firstIdx,
      cmd_lastIdx                              => s_read_first_name_cmd_lastIdx,
      cmd_ctrl                                 => s_read_first_name_cmd_ctrl,
      cmd_tag                                  => s_read_first_name_cmd_tag,
      unlock_valid                             => s_read_first_name_unlock_valid,
      unlock_ready                             => s_read_first_name_unlock_ready,
      unlock_tag                               => s_read_first_name_unlock_tag,
      out_valid                                => s_read_first_name_out_valid,
      out_ready                                => s_read_first_name_out_ready,
      out_last                                 => s_read_first_name_out_last,
      out_data                                 => s_read_first_name_out_data,
      out_dvalid                               => s_read_first_name_out_dvalid,
      bus_rreq_valid                           => s_read_first_name_bus_rreq_valid,
      bus_rreq_ready                           => s_read_first_name_bus_rreq_ready,
      bus_rreq_addr                            => s_read_first_name_bus_rreq_addr,
      bus_rreq_len                             => s_read_first_name_bus_rreq_len,
      bus_rdat_valid                           => s_read_first_name_bus_rdat_valid,
      bus_rdat_ready                           => s_read_first_name_bus_rdat_ready,
      bus_rdat_data                            => s_read_first_name_bus_rdat_data,
      bus_rdat_last                            => s_read_first_name_bus_rdat_last
    );

  -- ArrayReader instance generated from Arrow schema field:
  -- read_last_name: string not null
  read_last_name_read_inst: ArrayReader
    generic map (
      CFG                                      => "listprim(8)",
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH                            => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH                           => BUS_DATA_WIDTH,
      BUS_BURST_STEP_LEN                       => BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN                        => BUS_BURST_MAX_LEN,
      INDEX_WIDTH                              => INDEX_WIDTH,
      CMD_TAG_WIDTH                            => TAG_WIDTH,
      CMD_TAG_ENABLE                           => true
    )
    port map (
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      cmd_valid                                => s_read_last_name_cmd_valid,
      cmd_ready                                => s_read_last_name_cmd_ready,
      cmd_firstIdx                             => s_read_last_name_cmd_firstIdx,
      cmd_lastIdx                              => s_read_last_name_cmd_lastIdx,
      cmd_ctrl                                 => s_read_last_name_cmd_ctrl,
      cmd_tag                                  => s_read_last_name_cmd_tag,
      unlock_valid                             => s_read_last_name_unlock_valid,
      unlock_ready                             => s_read_last_name_unlock_ready,
      unlock_tag                               => s_read_last_name_unlock_tag,
      out_valid                                => s_read_last_name_out_valid,
      out_ready                                => s_read_last_name_out_ready,
      out_last                                 => s_read_last_name_out_last,
      out_data                                 => s_read_last_name_out_data,
      out_dvalid                               => s_read_last_name_out_dvalid,
      bus_rreq_valid                           => s_read_last_name_bus_rreq_valid,
      bus_rreq_ready                           => s_read_last_name_bus_rreq_ready,
      bus_rreq_addr                            => s_read_last_name_bus_rreq_addr,
      bus_rreq_len                             => s_read_last_name_bus_rreq_len,
      bus_rdat_valid                           => s_read_last_name_bus_rdat_valid,
      bus_rdat_ready                           => s_read_last_name_bus_rdat_ready,
      bus_rdat_data                            => s_read_last_name_bus_rdat_data,
      bus_rdat_last                            => s_read_last_name_bus_rdat_last
    );

  -- ArrayReader instance generated from Arrow schema field:
  -- read_zipcode: uint32 not null
  read_zipcode_read_inst: ArrayReader
    generic map (
      CFG                                      => "prim(32)",
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH                            => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH                           => BUS_DATA_WIDTH,
      BUS_BURST_STEP_LEN                       => BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN                        => BUS_BURST_MAX_LEN,
      INDEX_WIDTH                              => INDEX_WIDTH,
      CMD_TAG_WIDTH                            => TAG_WIDTH,
      CMD_TAG_ENABLE                           => true
    )
    port map (
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      cmd_valid                                => s_read_zipcode_cmd_valid,
      cmd_ready                                => s_read_zipcode_cmd_ready,
      cmd_firstIdx                             => s_read_zipcode_cmd_firstIdx,
      cmd_lastIdx                              => s_read_zipcode_cmd_lastIdx,
      cmd_ctrl                                 => s_read_zipcode_cmd_ctrl,
      cmd_tag                                  => s_read_zipcode_cmd_tag,
      unlock_valid                             => s_read_zipcode_unlock_valid,
      unlock_ready                             => s_read_zipcode_unlock_ready,
      unlock_tag                               => s_read_zipcode_unlock_tag,
      out_valid                                => s_read_zipcode_out_valid,
      out_ready                                => s_read_zipcode_out_ready,
      out_last                                 => s_read_zipcode_out_last,
      out_data                                 => s_read_zipcode_out_data,
      out_dvalid                               => s_read_zipcode_out_dvalid,
      bus_rreq_valid                           => s_read_zipcode_bus_rreq_valid,
      bus_rreq_ready                           => s_read_zipcode_bus_rreq_ready,
      bus_rreq_addr                            => s_read_zipcode_bus_rreq_addr,
      bus_rreq_len                             => s_read_zipcode_bus_rreq_len,
      bus_rdat_valid                           => s_read_zipcode_bus_rdat_valid,
      bus_rdat_ready                           => s_read_zipcode_bus_rdat_ready,
      bus_rdat_data                            => s_read_zipcode_bus_rdat_data,
      bus_rdat_last                            => s_read_zipcode_bus_rdat_last
    );

  -- ArrayWriter instance generated from Arrow schema field:
  -- write_first_name: string not null
  write_first_name_write_inst: ArrayWriter
    generic map (
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH                            => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH                           => BUS_DATA_WIDTH,
      BUS_STROBE_WIDTH                         => BUS_STROBE_WIDTH,
      BUS_BURST_STEP_LEN                       => BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN                        => BUS_BURST_MAX_LEN,
      INDEX_WIDTH                              => INDEX_WIDTH,
      CFG                                      => "listprim(8;last_from_length=0)",
      CMD_TAG_WIDTH                            => TAG_WIDTH,
      CMD_TAG_ENABLE                           => true
    )
    port map (
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      cmd_valid                                => s_write_first_name_cmd_valid,
      cmd_ready                                => s_write_first_name_cmd_ready,
      cmd_firstIdx                             => s_write_first_name_cmd_firstIdx,
      cmd_lastIdx                              => s_write_first_name_cmd_lastIdx,
      cmd_ctrl                                 => s_write_first_name_cmd_ctrl,
      cmd_tag                                  => s_write_first_name_cmd_tag,
      unlock_valid                             => s_write_first_name_unlock_valid,
      unlock_ready                             => s_write_first_name_unlock_ready,
      unlock_tag                               => s_write_first_name_unlock_tag,
      in_valid                                 => s_write_first_name_in_valid,
      in_ready                                 => s_write_first_name_in_ready,
      in_last                                  => s_write_first_name_in_last,
      in_data                                  => s_write_first_name_in_data,
      in_dvalid                                => s_write_first_name_in_dvalid,
      bus_wreq_valid                           => s_write_first_name_bus_wreq_valid,
      bus_wreq_ready                           => s_write_first_name_bus_wreq_ready,
      bus_wreq_addr                            => s_write_first_name_bus_wreq_addr,
      bus_wreq_len                             => s_write_first_name_bus_wreq_len,
      bus_wdat_valid                           => s_write_first_name_bus_wdat_valid,
      bus_wdat_ready                           => s_write_first_name_bus_wdat_ready,
      bus_wdat_data                            => s_write_first_name_bus_wdat_data,
      bus_wdat_strobe                          => s_write_first_name_bus_wdat_strobe,
      bus_wdat_last                            => s_write_first_name_bus_wdat_last
    );

  -- Controller instance.
  UserCoreController_inst: UserCoreController
    generic map (
      REG_WIDTH                                => REG_WIDTH
    )
    port map (
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      status                                   => regs_out(2*REG_WIDTH-1 downto REG_WIDTH),
      control                                  => regs_in(REG_WIDTH-1 downto 0),
      start                                    => uctrl_start,
      stop                                     => uctrl_stop,
      reset                                    => uctrl_reset,
      idle                                     => uctrl_idle,
      busy                                     => uctrl_busy,
      done                                     => uctrl_done
    );

  -- Hardware Accelerated Function instance.
  filter_usercore_inst: filter_usercore
    generic map (
      TAG_WIDTH                                => TAG_WIDTH,
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      INDEX_WIDTH                              => INDEX_WIDTH,
      REG_WIDTH                                => REG_WIDTH
    )
    port map (
      acc_clk                                  => acc_clk,
      acc_reset                                => acc_reset,
      ctrl_start                               => uctrl_start,
      ctrl_stop                                => uctrl_stop,
      ctrl_reset                               => uctrl_reset,
      ctrl_idle                                => uctrl_idle,
      ctrl_busy                                => uctrl_busy,
      ctrl_done                                => uctrl_done,
      read_first_name_out_valid                => s_read_first_name_out_valid(0),
      read_first_name_out_ready                => s_read_first_name_out_ready(0),
      read_first_name_out_last                 => s_read_first_name_out_last(0),
      read_first_name_out_length               => s_read_first_name_out_data(INDEX_WIDTH-1 downto 0),
      read_first_name_out_values_out_valid     => s_read_first_name_out_valid(1),
      read_first_name_out_values_out_ready     => s_read_first_name_out_ready(1),
      read_first_name_out_values_out_last      => s_read_first_name_out_last(1),
      read_first_name_out_values_out_dvalid    => s_read_first_name_out_dvalid(1),
      read_first_name_out_values_out_data      => s_read_first_name_out_data(INDEX_WIDTH+7 downto INDEX_WIDTH),
      read_first_name_out_values_out_count     => s_read_first_name_out_data(INDEX_WIDTH+8 downto INDEX_WIDTH+8),
      read_first_name_cmd_valid                => s_read_first_name_cmd_valid,
      read_first_name_cmd_ready                => s_read_first_name_cmd_ready,
      read_first_name_cmd_firstIdx             => s_read_first_name_cmd_firstIdx(INDEX_WIDTH-1 downto 0),
      read_first_name_cmd_lastIdx              => s_read_first_name_cmd_lastIdx(INDEX_WIDTH-1 downto 0),
      read_first_name_cmd_tag                  => s_read_first_name_cmd_tag(TAG_WIDTH-1 downto 0),
      read_first_name_cmd_read_first_name_offsets_addr=> s_read_first_name_cmd_ctrl(BUS_ADDR_WIDTH-1 downto 0),
      read_first_name_cmd_read_first_name_values_addr=> s_read_first_name_cmd_ctrl(BUS_ADDR_WIDTH+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH),
      read_first_name_unlock_valid             => s_read_first_name_unlock_valid,
      read_first_name_unlock_ready             => s_read_first_name_unlock_ready,
      read_first_name_unlock_tag               => s_read_first_name_unlock_tag,
      read_last_name_out_valid                 => s_read_last_name_out_valid(0),
      read_last_name_out_ready                 => s_read_last_name_out_ready(0),
      read_last_name_out_last                  => s_read_last_name_out_last(0),
      read_last_name_out_length                => s_read_last_name_out_data(INDEX_WIDTH-1 downto 0),
      read_last_name_out_values_out_valid      => s_read_last_name_out_valid(1),
      read_last_name_out_values_out_ready      => s_read_last_name_out_ready(1),
      read_last_name_out_values_out_last       => s_read_last_name_out_last(1),
      read_last_name_out_values_out_dvalid     => s_read_last_name_out_dvalid(1),
      read_last_name_out_values_out_data       => s_read_last_name_out_data(INDEX_WIDTH+7 downto INDEX_WIDTH),
      read_last_name_out_values_out_count      => s_read_last_name_out_data(INDEX_WIDTH+8 downto INDEX_WIDTH+8),
      read_last_name_cmd_valid                 => s_read_last_name_cmd_valid,
      read_last_name_cmd_ready                 => s_read_last_name_cmd_ready,
      read_last_name_cmd_firstIdx              => s_read_last_name_cmd_firstIdx(INDEX_WIDTH-1 downto 0),
      read_last_name_cmd_lastIdx               => s_read_last_name_cmd_lastIdx(INDEX_WIDTH-1 downto 0),
      read_last_name_cmd_tag                   => s_read_last_name_cmd_tag(TAG_WIDTH-1 downto 0),
      read_last_name_cmd_read_last_name_offsets_addr=> s_read_last_name_cmd_ctrl(BUS_ADDR_WIDTH-1 downto 0),
      read_last_name_cmd_read_last_name_values_addr=> s_read_last_name_cmd_ctrl(BUS_ADDR_WIDTH+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH),
      read_last_name_unlock_valid              => s_read_last_name_unlock_valid,
      read_last_name_unlock_ready              => s_read_last_name_unlock_ready,
      read_last_name_unlock_tag                => s_read_last_name_unlock_tag,
      read_zipcode_out_valid                   => s_read_zipcode_out_valid(0),
      read_zipcode_out_ready                   => s_read_zipcode_out_ready(0),
      read_zipcode_out_last                    => s_read_zipcode_out_last(0),
      read_zipcode_out_data                    => s_read_zipcode_out_data(31 downto 0),
      read_zipcode_cmd_valid                   => s_read_zipcode_cmd_valid,
      read_zipcode_cmd_ready                   => s_read_zipcode_cmd_ready,
      read_zipcode_cmd_firstIdx                => s_read_zipcode_cmd_firstIdx(INDEX_WIDTH-1 downto 0),
      read_zipcode_cmd_lastIdx                 => s_read_zipcode_cmd_lastIdx(INDEX_WIDTH-1 downto 0),
      read_zipcode_cmd_tag                     => s_read_zipcode_cmd_tag(TAG_WIDTH-1 downto 0),
      read_zipcode_cmd_read_zipcode_values_addr=> s_read_zipcode_cmd_ctrl(BUS_ADDR_WIDTH-1 downto 0),
      read_zipcode_unlock_valid                => s_read_zipcode_unlock_valid,
      read_zipcode_unlock_ready                => s_read_zipcode_unlock_ready,
      read_zipcode_unlock_tag                  => s_read_zipcode_unlock_tag,
      write_first_name_in_valid                => s_write_first_name_in_valid(0),
      write_first_name_in_ready                => s_write_first_name_in_ready(0),
      write_first_name_in_last                 => s_write_first_name_in_last(0),
      write_first_name_in_length               => s_write_first_name_in_data(INDEX_WIDTH-1 downto 0),
      write_first_name_in_values_in_valid      => s_write_first_name_in_valid(1),
      write_first_name_in_values_in_ready      => s_write_first_name_in_ready(1),
      write_first_name_in_values_in_last       => s_write_first_name_in_last(1),
      write_first_name_in_values_in_dvalid     => s_write_first_name_in_dvalid(1),
      write_first_name_in_values_in_data       => s_write_first_name_in_data(INDEX_WIDTH+7 downto INDEX_WIDTH),
      write_first_name_in_values_in_count      => s_write_first_name_in_data(INDEX_WIDTH+8 downto INDEX_WIDTH+8),
      write_first_name_cmd_valid               => s_write_first_name_cmd_valid,
      write_first_name_cmd_ready               => s_write_first_name_cmd_ready,
      write_first_name_cmd_firstIdx            => s_write_first_name_cmd_firstIdx(INDEX_WIDTH-1 downto 0),
      write_first_name_cmd_lastIdx             => s_write_first_name_cmd_lastIdx(INDEX_WIDTH-1 downto 0),
      write_first_name_cmd_tag                 => s_write_first_name_cmd_tag(TAG_WIDTH-1 downto 0),
      write_first_name_cmd_write_first_name_offsets_addr=> s_write_first_name_cmd_ctrl(BUS_ADDR_WIDTH-1 downto 0),
      write_first_name_cmd_write_first_name_values_addr=> s_write_first_name_cmd_ctrl(BUS_ADDR_WIDTH+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH),
      write_first_name_unlock_valid            => s_write_first_name_unlock_valid,
      write_first_name_unlock_ready            => s_write_first_name_unlock_ready,
      write_first_name_unlock_tag              => s_write_first_name_unlock_tag,
      idx_first                                => regs_in(5*REG_WIDTH-1 downto 4*REG_WIDTH),
      idx_last                                 => regs_in(6*REG_WIDTH-1 downto 5*REG_WIDTH),
      reg_return0                              => regs_out(3*REG_WIDTH-1 downto 2*REG_WIDTH),
      reg_return1                              => regs_out(4*REG_WIDTH-1 downto 3*REG_WIDTH),
      reg_read_first_name_offsets_addr         => regs_in(8*REG_WIDTH-1 downto 6*REG_WIDTH),
      reg_read_first_name_values_addr          => regs_in(10*REG_WIDTH-1 downto 8*REG_WIDTH),
      reg_read_last_name_offsets_addr          => regs_in(12*REG_WIDTH-1 downto 10*REG_WIDTH),
      reg_read_last_name_values_addr           => regs_in(14*REG_WIDTH-1 downto 12*REG_WIDTH),
      reg_read_zipcode_values_addr             => regs_in(16*REG_WIDTH-1 downto 14*REG_WIDTH),
      reg_write_first_name_offsets_addr        => regs_in(18*REG_WIDTH-1 downto 16*REG_WIDTH),
      reg_write_first_name_values_addr         => regs_in(20*REG_WIDTH-1 downto 18*REG_WIDTH)
    );

  -- Arbiter instance generated to serve 3 array readers.
  BusReadArbiterVec_inst: BusReadArbiterVec
    generic map (
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH                            => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH                           => BUS_DATA_WIDTH,
      NUM_SLAVE_PORTS                          => 3
    )
    port map (
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      bsv_rreq_valid                           => s_bsv_rreq_valid,
      bsv_rreq_ready                           => s_bsv_rreq_ready,
      bsv_rreq_addr                            => s_bsv_rreq_addr,
      bsv_rreq_len                             => s_bsv_rreq_len,
      bsv_rdat_valid                           => s_bsv_rdat_valid,
      bsv_rdat_ready                           => s_bsv_rdat_ready,
      bsv_rdat_data                            => s_bsv_rdat_data,
      bsv_rdat_last                            => s_bsv_rdat_last,
      mst_rreq_valid                           => mst_rreq_valid,
      mst_rreq_ready                           => mst_rreq_ready,
      mst_rreq_addr                            => mst_rreq_addr,
      mst_rreq_len                             => mst_rreq_len,
      mst_rdat_valid                           => mst_rdat_valid,
      mst_rdat_ready                           => mst_rdat_ready,
      mst_rdat_data                            => mst_rdat_data,
      mst_rdat_last                            => mst_rdat_last
    );

  -- Arbiter instance generated to serve 1 array writers.
  BusWriteArbiterVec_inst: BusWriteArbiterVec
    generic map (
      BUS_ADDR_WIDTH                           => BUS_ADDR_WIDTH,
      BUS_LEN_WIDTH                            => BUS_LEN_WIDTH,
      BUS_DATA_WIDTH                           => BUS_DATA_WIDTH,
      BUS_STROBE_WIDTH                         => BUS_STROBE_WIDTH,
      NUM_SLAVE_PORTS                          => 1
    )
    port map (
      bus_clk                                  => bus_clk,
      bus_reset                                => bus_reset,
      bsv_wdat_valid                           => s_bsv_wdat_valid,
      bsv_wdat_ready                           => s_bsv_wdat_ready,
      bsv_wdat_data                            => s_bsv_wdat_data,
      bsv_wdat_strobe                          => s_bsv_wdat_strobe,
      bsv_wdat_last                            => s_bsv_wdat_last,
      bsv_wreq_valid                           => s_bsv_wreq_valid,
      bsv_wreq_ready                           => s_bsv_wreq_ready,
      bsv_wreq_addr                            => s_bsv_wreq_addr,
      bsv_wreq_len                             => s_bsv_wreq_len,
      mst_wreq_valid                           => mst_wreq_valid,
      mst_wreq_ready                           => mst_wreq_ready,
      mst_wreq_addr                            => mst_wreq_addr,
      mst_wreq_len                             => mst_wreq_len,
      mst_wdat_valid                           => mst_wdat_valid,
      mst_wdat_ready                           => mst_wdat_ready,
      mst_wdat_data                            => mst_wdat_data,
      mst_wdat_strobe                          => mst_wdat_strobe,
      mst_wdat_last                            => mst_wdat_last
    );


  s_bsv_rreq_valid(0)                          <= s_read_first_name_bus_rreq_valid;
  s_read_first_name_bus_rreq_ready             <= s_bsv_rreq_ready(0);
  s_bsv_rreq_len(BUS_LEN_WIDTH-1 downto 0)     <= s_read_first_name_bus_rreq_len;
  s_bsv_rreq_addr(BUS_ADDR_WIDTH-1 downto 0)   <= s_read_first_name_bus_rreq_addr;
  -----------------------------------------------------------------------------
  s_bsv_rreq_valid(1)                          <= s_read_last_name_bus_rreq_valid;
  s_read_last_name_bus_rreq_ready              <= s_bsv_rreq_ready(1);
  s_bsv_rreq_len(2*BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH)<= s_read_last_name_bus_rreq_len;
  s_bsv_rreq_addr(2*BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH)<= s_read_last_name_bus_rreq_addr;
  -----------------------------------------------------------------------------
  s_bsv_rreq_valid(2)                          <= s_read_zipcode_bus_rreq_valid;
  s_read_zipcode_bus_rreq_ready                <= s_bsv_rreq_ready(2);
  s_bsv_rreq_len(3*BUS_LEN_WIDTH-1 downto 2*BUS_LEN_WIDTH)<= s_read_zipcode_bus_rreq_len;
  s_bsv_rreq_addr(3*BUS_ADDR_WIDTH-1 downto 2*BUS_ADDR_WIDTH)<= s_read_zipcode_bus_rreq_addr;
  -----------------------------------------------------------------------------
  s_read_first_name_bus_rdat_data              <= s_bsv_rdat_data(BUS_DATA_WIDTH-1 downto 0);
  s_read_first_name_bus_rdat_valid             <= s_bsv_rdat_valid(0);
  s_bsv_rdat_ready(0)                          <= s_read_first_name_bus_rdat_ready;
  s_read_first_name_bus_rdat_last              <= s_bsv_rdat_last(0);
  -----------------------------------------------------------------------------
  s_read_last_name_bus_rdat_data               <= s_bsv_rdat_data(2*BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH);
  s_read_last_name_bus_rdat_valid              <= s_bsv_rdat_valid(1);
  s_read_last_name_bus_rdat_last               <= s_bsv_rdat_last(1);
  s_bsv_rdat_ready(1)                          <= s_read_last_name_bus_rdat_ready;
  -----------------------------------------------------------------------------
  s_read_zipcode_bus_rdat_last                 <= s_bsv_rdat_last(2);
  s_bsv_rdat_ready(2)                          <= s_read_zipcode_bus_rdat_ready;
  s_read_zipcode_bus_rdat_data                 <= s_bsv_rdat_data(3*BUS_DATA_WIDTH-1 downto 2*BUS_DATA_WIDTH);
  s_read_zipcode_bus_rdat_valid                <= s_bsv_rdat_valid(2);
  -----------------------------------------------------------------------------
  s_bsv_wreq_addr(BUS_ADDR_WIDTH-1 downto 0)   <= s_write_first_name_bus_wreq_addr;
  s_bsv_wreq_len(BUS_LEN_WIDTH-1 downto 0)     <= s_write_first_name_bus_wreq_len;
  s_write_first_name_bus_wreq_ready            <= s_bsv_wreq_ready(0);
  s_bsv_wreq_valid(0)                          <= s_write_first_name_bus_wreq_valid;
  -----------------------------------------------------------------------------
  s_bsv_wdat_data(BUS_DATA_WIDTH-1 downto 0)   <= s_write_first_name_bus_wdat_data;
  s_bsv_wdat_last(0)                           <= s_write_first_name_bus_wdat_last;
  s_write_first_name_bus_wdat_ready            <= s_bsv_wdat_ready(0);
  s_bsv_wdat_strobe(BUS_STROBE_WIDTH-1 downto 0)<= s_write_first_name_bus_wdat_strobe;
  s_bsv_wdat_valid(0)                          <= s_write_first_name_bus_wdat_valid;
  -----------------------------------------------------------------------------
  regs_out_en(0)                               <='0';
  regs_out_en(1)                               <='1';
  regs_out_en(2)                               <='1';
  regs_out_en(3)                               <='1';

end architecture;

